VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 87.460 2924.800 88.660 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2433.460 2924.800 2434.660 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 2866.000 2663.660 2901.150 2663.800 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
      LAYER via ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
      LAYER met2 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
      LAYER met3 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 2866.000 2898.260 2901.150 2898.400 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
      LAYER via ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 2866.000 3132.860 2901.150 3133.000 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
      LAYER via ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 2866.000 3367.460 2901.150 3367.600 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
      LAYER via ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2445.890 3501.560 2446.210 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 2445.890 3501.420 2798.570 3501.560 ;
        RECT 2445.890 3501.360 2446.210 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
      LAYER via ;
        RECT 2445.920 3501.360 2446.180 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 2445.920 3501.330 2446.180 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 2445.980 3466.000 2446.120 3501.330 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2452.790 3498.500 2453.110 3498.560 ;
        RECT 2473.950 3498.500 2474.270 3498.560 ;
        RECT 2452.790 3498.360 2474.270 3498.500 ;
        RECT 2452.790 3498.300 2453.110 3498.360 ;
        RECT 2473.950 3498.300 2474.270 3498.360 ;
      LAYER via ;
        RECT 2452.820 3498.300 2453.080 3498.560 ;
        RECT 2473.980 3498.300 2474.240 3498.560 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3498.590 2474.180 3517.600 ;
        RECT 2452.820 3498.270 2453.080 3498.590 ;
        RECT 2473.980 3498.270 2474.240 3498.590 ;
        RECT 2452.880 3466.000 2453.020 3498.270 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2149.190 3498.500 2149.510 3498.560 ;
        RECT 2152.410 3498.500 2152.730 3498.560 ;
        RECT 2149.190 3498.360 2152.730 3498.500 ;
        RECT 2149.190 3498.300 2149.510 3498.360 ;
        RECT 2152.410 3498.300 2152.730 3498.360 ;
      LAYER via ;
        RECT 2149.220 3498.300 2149.480 3498.560 ;
        RECT 2152.440 3498.300 2152.700 3498.560 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3498.590 2149.420 3517.600 ;
        RECT 2149.220 3498.270 2149.480 3498.590 ;
        RECT 2152.440 3498.270 2152.700 3498.590 ;
        RECT 2152.500 3466.000 2152.640 3498.270 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1824.890 3498.500 1825.210 3498.560 ;
        RECT 1828.110 3498.500 1828.430 3498.560 ;
        RECT 1824.890 3498.360 1828.430 3498.500 ;
        RECT 1824.890 3498.300 1825.210 3498.360 ;
        RECT 1828.110 3498.300 1828.430 3498.360 ;
      LAYER via ;
        RECT 1824.920 3498.300 1825.180 3498.560 ;
        RECT 1828.140 3498.300 1828.400 3498.560 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3498.590 1825.120 3517.600 ;
        RECT 1824.920 3498.270 1825.180 3498.590 ;
        RECT 1828.140 3498.270 1828.400 3498.590 ;
        RECT 1828.200 3466.000 1828.340 3498.270 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3498.500 1500.910 3498.560 ;
        RECT 1503.810 3498.500 1504.130 3498.560 ;
        RECT 1500.590 3498.360 1504.130 3498.500 ;
        RECT 1500.590 3498.300 1500.910 3498.360 ;
        RECT 1503.810 3498.300 1504.130 3498.360 ;
      LAYER via ;
        RECT 1500.620 3498.300 1500.880 3498.560 ;
        RECT 1503.840 3498.300 1504.100 3498.560 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3498.590 1500.820 3517.600 ;
        RECT 1500.620 3498.270 1500.880 3498.590 ;
        RECT 1503.840 3498.270 1504.100 3498.590 ;
        RECT 1503.900 3466.000 1504.040 3498.270 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 322.060 2924.800 323.260 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 3466.000 1179.740 3498.270 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3498.500 851.850 3498.560 ;
        RECT 855.210 3498.500 855.530 3498.560 ;
        RECT 851.530 3498.360 855.530 3498.500 ;
        RECT 851.530 3498.300 851.850 3498.360 ;
        RECT 855.210 3498.300 855.530 3498.360 ;
      LAYER via ;
        RECT 851.560 3498.300 851.820 3498.560 ;
        RECT 855.240 3498.300 855.500 3498.560 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3498.590 851.760 3517.600 ;
        RECT 851.560 3498.270 851.820 3498.590 ;
        RECT 855.240 3498.270 855.500 3498.590 ;
        RECT 855.300 3466.000 855.440 3498.270 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.910 3498.500 531.230 3498.560 ;
        RECT 527.230 3498.360 531.230 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.910 3498.300 531.230 3498.360 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.940 3498.300 531.200 3498.560 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.940 3498.270 531.200 3498.590 ;
        RECT 531.000 3466.000 531.140 3498.270 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3502.580 202.790 3502.640 ;
        RECT 206.610 3502.580 206.930 3502.640 ;
        RECT 202.470 3502.440 206.930 3502.580 ;
        RECT 202.470 3502.380 202.790 3502.440 ;
        RECT 206.610 3502.380 206.930 3502.440 ;
      LAYER via ;
        RECT 202.500 3502.380 202.760 3502.640 ;
        RECT 206.640 3502.380 206.900 3502.640 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3502.670 202.700 3517.600 ;
        RECT 202.500 3502.350 202.760 3502.670 ;
        RECT 206.640 3502.350 206.900 3502.670 ;
        RECT 206.700 3466.000 206.840 3502.350 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 17.550 3408.600 54.000 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 3119.060 17.410 3119.120 ;
        RECT 17.090 3118.920 54.000 3119.060 ;
        RECT 17.090 3118.860 17.410 3118.920 ;
      LAYER via ;
        RECT 17.120 3118.860 17.380 3119.120 ;
      LAYER met2 ;
        RECT 17.110 3124.075 17.390 3124.445 ;
        RECT 17.180 3119.150 17.320 3124.075 ;
        RECT 17.120 3118.830 17.380 3119.150 ;
      LAYER via2 ;
        RECT 17.110 3124.120 17.390 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.085 3124.410 17.415 3124.425 ;
        RECT -4.800 3124.110 17.415 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.085 3124.095 17.415 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2836.180 17.410 2836.240 ;
        RECT 17.090 2836.040 54.000 2836.180 ;
        RECT 17.090 2835.980 17.410 2836.040 ;
      LAYER via ;
        RECT 17.120 2835.980 17.380 2836.240 ;
      LAYER met2 ;
        RECT 17.110 2836.435 17.390 2836.805 ;
        RECT 17.180 2836.270 17.320 2836.435 ;
        RECT 17.120 2835.950 17.380 2836.270 ;
      LAYER via2 ;
        RECT 17.110 2836.480 17.390 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 17.085 2836.770 17.415 2836.785 ;
        RECT -4.800 2836.470 17.415 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 17.085 2836.455 17.415 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2549.060 2.400 2550.260 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2261.420 2.400 2262.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1974.460 2.400 1975.660 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 556.660 2924.800 557.860 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1686.820 2.400 1688.020 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1471.260 2.400 1472.460 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1255.700 2.400 1256.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1040.140 2.400 1041.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 824.580 2.400 825.780 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 609.700 2.400 610.900 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 394.140 2.400 395.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 178.580 2.400 179.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 791.260 2924.800 792.460 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1025.860 2924.800 1027.060 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1260.460 2924.800 1261.660 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1495.060 2924.800 1496.260 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1729.660 2924.800 1730.860 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1964.260 2924.800 1965.460 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2198.860 2924.800 2200.060 ;
    END
  END io_in[9]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 2866.000 2780.960 2901.150 2781.100 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
      LAYER via ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 2866.000 3015.560 2901.150 3015.700 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 2866.000 3250.160 2901.150 3250.300 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
      LAYER via ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2480.390 3484.900 2480.710 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 2480.390 3484.760 2901.150 3484.900 ;
        RECT 2480.390 3484.700 2480.710 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 2480.420 3484.700 2480.680 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 2480.420 3484.670 2480.680 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 2480.480 3466.000 2480.620 3484.670 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2487.290 3502.240 2487.610 3502.300 ;
        RECT 2635.870 3502.240 2636.190 3502.300 ;
        RECT 2487.290 3502.100 2636.190 3502.240 ;
        RECT 2487.290 3502.040 2487.610 3502.100 ;
        RECT 2635.870 3502.040 2636.190 3502.100 ;
      LAYER via ;
        RECT 2487.320 3502.040 2487.580 3502.300 ;
        RECT 2635.900 3502.040 2636.160 3502.300 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3502.330 2636.100 3517.600 ;
        RECT 2487.320 3502.010 2487.580 3502.330 ;
        RECT 2635.900 3502.010 2636.160 3502.330 ;
        RECT 2487.380 3466.000 2487.520 3502.010 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2311.570 3498.500 2311.890 3498.560 ;
        RECT 2318.010 3498.500 2318.330 3498.560 ;
        RECT 2311.570 3498.360 2318.330 3498.500 ;
        RECT 2311.570 3498.300 2311.890 3498.360 ;
        RECT 2318.010 3498.300 2318.330 3498.360 ;
      LAYER via ;
        RECT 2311.600 3498.300 2311.860 3498.560 ;
        RECT 2318.040 3498.300 2318.300 3498.560 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3498.590 2311.800 3517.600 ;
        RECT 2311.600 3498.270 2311.860 3498.590 ;
        RECT 2318.040 3498.270 2318.300 3498.590 ;
        RECT 2318.100 3466.000 2318.240 3498.270 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1987.270 3499.860 1987.590 3499.920 ;
        RECT 1993.710 3499.860 1994.030 3499.920 ;
        RECT 1987.270 3499.720 1994.030 3499.860 ;
        RECT 1987.270 3499.660 1987.590 3499.720 ;
        RECT 1993.710 3499.660 1994.030 3499.720 ;
      LAYER via ;
        RECT 1987.300 3499.660 1987.560 3499.920 ;
        RECT 1993.740 3499.660 1994.000 3499.920 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3499.950 1987.500 3517.600 ;
        RECT 1987.300 3499.630 1987.560 3499.950 ;
        RECT 1993.740 3499.630 1994.000 3499.950 ;
        RECT 1993.800 3466.000 1993.940 3499.630 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3466.000 1662.740 3517.600 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3503.600 1338.530 3503.660 ;
        RECT 2401.270 3503.600 2401.590 3503.660 ;
        RECT 1338.210 3503.460 2401.590 3503.600 ;
        RECT 1338.210 3503.400 1338.530 3503.460 ;
        RECT 2401.270 3503.400 2401.590 3503.460 ;
      LAYER via ;
        RECT 1338.240 3503.400 1338.500 3503.660 ;
        RECT 2401.300 3503.400 2401.560 3503.660 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3503.690 1338.440 3517.600 ;
        RECT 1338.240 3503.370 1338.500 3503.690 ;
        RECT 2401.300 3503.370 2401.560 3503.690 ;
        RECT 2401.360 3466.000 2401.500 3503.370 ;
    END
  END io_oeb[19]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3503.260 1014.230 3503.320 ;
        RECT 2391.150 3503.260 2391.470 3503.320 ;
        RECT 1013.910 3503.120 2391.470 3503.260 ;
        RECT 1013.910 3503.060 1014.230 3503.120 ;
        RECT 2391.150 3503.060 2391.470 3503.120 ;
      LAYER via ;
        RECT 1013.940 3503.060 1014.200 3503.320 ;
        RECT 2391.180 3503.060 2391.440 3503.320 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3503.350 1014.140 3517.600 ;
        RECT 1013.940 3503.030 1014.200 3503.350 ;
        RECT 2391.180 3503.030 2391.440 3503.350 ;
        RECT 2391.240 3466.000 2391.380 3503.030 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3502.920 689.470 3502.980 ;
        RECT 2391.610 3502.920 2391.930 3502.980 ;
        RECT 689.150 3502.780 2391.930 3502.920 ;
        RECT 689.150 3502.720 689.470 3502.780 ;
        RECT 2391.610 3502.720 2391.930 3502.780 ;
      LAYER via ;
        RECT 689.180 3502.720 689.440 3502.980 ;
        RECT 2391.640 3502.720 2391.900 3502.980 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3503.010 689.380 3517.600 ;
        RECT 689.180 3502.690 689.440 3503.010 ;
        RECT 2391.640 3502.690 2391.900 3503.010 ;
        RECT 2391.700 3466.000 2391.840 3502.690 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 3502.240 365.170 3502.300 ;
        RECT 2392.070 3502.240 2392.390 3502.300 ;
        RECT 364.850 3502.100 2392.390 3502.240 ;
        RECT 364.850 3502.040 365.170 3502.100 ;
        RECT 2392.070 3502.040 2392.390 3502.100 ;
      LAYER via ;
        RECT 364.880 3502.040 365.140 3502.300 ;
        RECT 2392.100 3502.040 2392.360 3502.300 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3502.330 365.080 3517.600 ;
        RECT 364.880 3502.010 365.140 3502.330 ;
        RECT 2392.100 3502.010 2392.360 3502.330 ;
        RECT 2392.160 3466.000 2392.300 3502.010 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.550 3501.560 40.870 3501.620 ;
        RECT 2387.470 3501.560 2387.790 3501.620 ;
        RECT 40.550 3501.420 2387.790 3501.560 ;
        RECT 40.550 3501.360 40.870 3501.420 ;
        RECT 2387.470 3501.360 2387.790 3501.420 ;
        RECT 2387.470 3498.500 2387.790 3498.560 ;
        RECT 2392.990 3498.500 2393.310 3498.560 ;
        RECT 2387.470 3498.360 2393.310 3498.500 ;
        RECT 2387.470 3498.300 2387.790 3498.360 ;
        RECT 2392.990 3498.300 2393.310 3498.360 ;
      LAYER via ;
        RECT 40.580 3501.360 40.840 3501.620 ;
        RECT 2387.500 3501.360 2387.760 3501.620 ;
        RECT 2387.500 3498.300 2387.760 3498.560 ;
        RECT 2393.020 3498.300 2393.280 3498.560 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.650 40.780 3517.600 ;
        RECT 40.580 3501.330 40.840 3501.650 ;
        RECT 2387.500 3501.330 2387.760 3501.650 ;
        RECT 2387.560 3498.590 2387.700 3501.330 ;
        RECT 2387.500 3498.270 2387.760 3498.590 ;
        RECT 2393.020 3498.270 2393.280 3498.590 ;
        RECT 2393.080 3466.000 2393.220 3498.270 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 15.250 3263.760 54.000 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 2974.220 16.490 2974.280 ;
        RECT 16.170 2974.080 54.000 2974.220 ;
        RECT 16.170 2974.020 16.490 2974.080 ;
      LAYER via ;
        RECT 16.200 2974.020 16.460 2974.280 ;
      LAYER met2 ;
        RECT 16.190 2979.915 16.470 2980.285 ;
        RECT 16.260 2974.310 16.400 2979.915 ;
        RECT 16.200 2973.990 16.460 2974.310 ;
      LAYER via2 ;
        RECT 16.190 2979.960 16.470 2980.240 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.165 2980.250 16.495 2980.265 ;
        RECT -4.800 2979.950 16.495 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.165 2979.935 16.495 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2691.340 17.410 2691.400 ;
        RECT 17.090 2691.200 54.000 2691.340 ;
        RECT 17.090 2691.140 17.410 2691.200 ;
      LAYER via ;
        RECT 17.120 2691.140 17.380 2691.400 ;
      LAYER met2 ;
        RECT 17.110 2692.955 17.390 2693.325 ;
        RECT 17.180 2691.430 17.320 2692.955 ;
        RECT 17.120 2691.110 17.380 2691.430 ;
      LAYER via2 ;
        RECT 17.110 2693.000 17.390 2693.280 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 17.085 2693.290 17.415 2693.305 ;
        RECT -4.800 2692.990 17.415 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 17.085 2692.975 17.415 2692.990 ;
    END
  END io_oeb[26]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 2866.000 2725.540 2901.150 2725.680 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
      LAYER via ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
      LAYER met3 ;
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 2866.000 2960.140 2901.150 2960.280 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
      LAYER via ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 2866.000 3194.740 2901.150 3194.880 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
      LAYER via ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2866.000 3429.340 2901.150 3429.480 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2521.790 3501.900 2522.110 3501.960 ;
        RECT 2717.290 3501.900 2717.610 3501.960 ;
        RECT 2521.790 3501.760 2717.610 3501.900 ;
        RECT 2521.790 3501.700 2522.110 3501.760 ;
        RECT 2717.290 3501.700 2717.610 3501.760 ;
      LAYER via ;
        RECT 2521.820 3501.700 2522.080 3501.960 ;
        RECT 2717.320 3501.700 2717.580 3501.960 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.990 2717.520 3517.600 ;
        RECT 2521.820 3501.670 2522.080 3501.990 ;
        RECT 2717.320 3501.670 2717.580 3501.990 ;
        RECT 2521.880 3466.000 2522.020 3501.670 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3499.010 2392.760 3517.600 ;
        RECT 2392.620 3498.870 2394.600 3499.010 ;
        RECT 2394.460 3466.000 2394.600 3498.870 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2068.230 3504.280 2068.550 3504.340 ;
        RECT 2389.770 3504.280 2390.090 3504.340 ;
        RECT 2068.230 3504.140 2390.090 3504.280 ;
        RECT 2068.230 3504.080 2068.550 3504.140 ;
        RECT 2389.770 3504.080 2390.090 3504.140 ;
      LAYER via ;
        RECT 2068.260 3504.080 2068.520 3504.340 ;
        RECT 2389.800 3504.080 2390.060 3504.340 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3504.370 2068.460 3517.600 ;
        RECT 2068.260 3504.050 2068.520 3504.370 ;
        RECT 2389.800 3504.050 2390.060 3504.370 ;
        RECT 2389.860 3497.650 2390.000 3504.050 ;
        RECT 2389.860 3497.510 2390.920 3497.650 ;
        RECT 2390.780 3466.000 2390.920 3497.510 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1743.930 3503.940 1744.250 3504.000 ;
        RECT 2394.830 3503.940 2395.150 3504.000 ;
        RECT 1743.930 3503.800 2395.150 3503.940 ;
        RECT 1743.930 3503.740 1744.250 3503.800 ;
        RECT 2394.830 3503.740 2395.150 3503.800 ;
      LAYER via ;
        RECT 1743.960 3503.740 1744.220 3504.000 ;
        RECT 2394.860 3503.740 2395.120 3504.000 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3504.030 1744.160 3517.600 ;
        RECT 1743.960 3503.710 1744.220 3504.030 ;
        RECT 2394.860 3503.710 2395.120 3504.030 ;
        RECT 2394.920 3466.000 2395.060 3503.710 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.170 3477.760 1419.490 3477.820 ;
        RECT 1419.630 3477.760 1419.950 3477.820 ;
        RECT 1419.170 3477.620 1419.950 3477.760 ;
        RECT 1419.170 3477.560 1419.490 3477.620 ;
        RECT 1419.630 3477.560 1419.950 3477.620 ;
      LAYER via ;
        RECT 1419.200 3477.560 1419.460 3477.820 ;
        RECT 1419.660 3477.560 1419.920 3477.820 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3477.850 1419.400 3517.600 ;
        RECT 1419.200 3477.530 1419.460 3477.850 ;
        RECT 1419.660 3477.530 1419.920 3477.850 ;
        RECT 1419.720 3466.000 1419.860 3477.530 ;
    END
  END io_out[19]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1095.405 3466.000 1095.575 3477.435 ;
      LAYER L1M1_PR_C ;
        RECT 1095.405 3477.265 1095.575 3477.435 ;
      LAYER met1 ;
        RECT 1095.345 3477.420 1095.635 3477.465 ;
        RECT 1095.790 3477.420 1096.110 3477.480 ;
        RECT 1095.345 3477.280 1096.110 3477.420 ;
        RECT 1095.345 3477.235 1095.635 3477.280 ;
        RECT 1095.790 3477.220 1096.110 3477.280 ;
      LAYER via ;
        RECT 1095.820 3477.220 1096.080 3477.480 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3517.370 1095.100 3517.600 ;
        RECT 1094.500 3517.230 1095.100 3517.370 ;
        RECT 1094.500 3478.725 1094.640 3517.230 ;
        RECT 1094.430 3478.355 1094.710 3478.725 ;
        RECT 1096.270 3477.930 1096.550 3478.045 ;
        RECT 1095.880 3477.790 1096.550 3477.930 ;
        RECT 1095.880 3477.510 1096.020 3477.790 ;
        RECT 1096.270 3477.675 1096.550 3477.790 ;
        RECT 1095.820 3477.190 1096.080 3477.510 ;
      LAYER via2 ;
        RECT 1094.430 3478.400 1094.710 3478.680 ;
        RECT 1096.270 3477.720 1096.550 3478.000 ;
      LAYER met3 ;
        RECT 1094.405 3478.690 1094.735 3478.705 ;
        RECT 1094.405 3478.390 1097.250 3478.690 ;
        RECT 1094.405 3478.375 1094.735 3478.390 ;
        RECT 1096.245 3478.010 1096.575 3478.025 ;
        RECT 1096.950 3478.010 1097.250 3478.390 ;
        RECT 1096.245 3477.710 1097.250 3478.010 ;
        RECT 1096.245 3477.695 1096.575 3477.710 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 770.570 3477.760 770.890 3477.820 ;
        RECT 771.030 3477.760 771.350 3477.820 ;
        RECT 770.570 3477.620 771.350 3477.760 ;
        RECT 770.570 3477.560 770.890 3477.620 ;
        RECT 771.030 3477.560 771.350 3477.620 ;
      LAYER via ;
        RECT 770.600 3477.560 770.860 3477.820 ;
        RECT 771.060 3477.560 771.320 3477.820 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3477.850 770.800 3517.600 ;
        RECT 770.600 3477.530 770.860 3477.850 ;
        RECT 771.060 3477.530 771.320 3477.850 ;
        RECT 771.120 3466.000 771.260 3477.530 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3502.580 446.130 3502.640 ;
        RECT 2390.690 3502.580 2391.010 3502.640 ;
        RECT 445.810 3502.440 2391.010 3502.580 ;
        RECT 445.810 3502.380 446.130 3502.440 ;
        RECT 2390.690 3502.380 2391.010 3502.440 ;
        RECT 2390.690 3498.160 2391.010 3498.220 ;
        RECT 2392.530 3498.160 2392.850 3498.220 ;
        RECT 2390.690 3498.020 2392.850 3498.160 ;
        RECT 2390.690 3497.960 2391.010 3498.020 ;
        RECT 2392.530 3497.960 2392.850 3498.020 ;
      LAYER via ;
        RECT 445.840 3502.380 446.100 3502.640 ;
        RECT 2390.720 3502.380 2390.980 3502.640 ;
        RECT 2390.720 3497.960 2390.980 3498.220 ;
        RECT 2392.560 3497.960 2392.820 3498.220 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3502.670 446.040 3517.600 ;
        RECT 445.840 3502.350 446.100 3502.670 ;
        RECT 2390.720 3502.350 2390.980 3502.670 ;
        RECT 2390.780 3498.250 2390.920 3502.350 ;
        RECT 2390.720 3497.930 2390.980 3498.250 ;
        RECT 2392.560 3497.930 2392.820 3498.250 ;
        RECT 2392.620 3466.000 2392.760 3497.930 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3501.900 121.830 3501.960 ;
        RECT 2395.290 3501.900 2395.610 3501.960 ;
        RECT 121.510 3501.760 2395.610 3501.900 ;
        RECT 121.510 3501.700 121.830 3501.760 ;
        RECT 2395.290 3501.700 2395.610 3501.760 ;
      LAYER via ;
        RECT 121.540 3501.700 121.800 3501.960 ;
        RECT 2395.320 3501.700 2395.580 3501.960 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3501.990 121.740 3517.600 ;
        RECT 121.540 3501.670 121.800 3501.990 ;
        RECT 2395.320 3501.670 2395.580 3501.990 ;
        RECT 2395.380 3466.000 2395.520 3501.670 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 17.090 3339.580 54.000 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3050.040 17.410 3050.100 ;
        RECT 17.090 3049.900 54.000 3050.040 ;
        RECT 17.090 3049.840 17.410 3049.900 ;
      LAYER via ;
        RECT 17.120 3049.840 17.380 3050.100 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3050.130 17.320 3051.995 ;
        RECT 17.120 3049.810 17.380 3050.130 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2760.360 16.030 2760.420 ;
        RECT 15.710 2760.220 54.000 2760.360 ;
        RECT 15.710 2760.160 16.030 2760.220 ;
      LAYER via ;
        RECT 15.740 2760.160 16.000 2760.420 ;
      LAYER met2 ;
        RECT 15.730 2765.035 16.010 2765.405 ;
        RECT 15.800 2760.450 15.940 2765.035 ;
        RECT 15.740 2760.130 16.000 2760.450 ;
      LAYER via2 ;
        RECT 15.730 2765.080 16.010 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 15.705 2765.370 16.035 2765.385 ;
        RECT -4.800 2765.070 16.035 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 15.705 2765.055 16.035 2765.070 ;
    END
  END io_out[26]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 48.445 1691.245 48.615 1692.435 ;
      LAYER L1M1_PR_C ;
        RECT 48.445 1692.265 48.615 1692.435 ;
      LAYER met1 ;
        RECT 48.385 1692.420 48.675 1692.465 ;
        RECT 48.385 1692.280 54.000 1692.420 ;
        RECT 48.385 1692.235 48.675 1692.280 ;
        RECT 17.090 1691.400 17.410 1691.460 ;
        RECT 48.385 1691.400 48.675 1691.445 ;
        RECT 17.090 1691.260 48.675 1691.400 ;
        RECT 17.090 1691.200 17.410 1691.260 ;
        RECT 48.385 1691.215 48.675 1691.260 ;
        RECT 2901.290 1690.720 2901.610 1690.780 ;
        RECT 2866.000 1690.580 2901.610 1690.720 ;
        RECT 2901.290 1690.520 2901.610 1690.580 ;
      LAYER via ;
        RECT 17.120 1691.200 17.380 1691.460 ;
        RECT 2901.320 1690.520 2901.580 1690.780 ;
      LAYER met2 ;
        RECT 2904.530 2551.515 2904.810 2551.885 ;
        RECT 2904.600 2493.405 2904.740 2551.515 ;
        RECT 2904.530 2493.035 2904.810 2493.405 ;
        RECT 13.890 2477.395 14.170 2477.765 ;
        RECT 13.960 2405.685 14.100 2477.395 ;
        RECT 13.890 2405.315 14.170 2405.685 ;
        RECT 13.960 2190.125 14.100 2405.315 ;
        RECT 2904.600 2317.285 2904.740 2493.035 ;
        RECT 2904.530 2316.915 2904.810 2317.285 ;
        RECT 2904.600 2258.805 2904.740 2316.915 ;
        RECT 2904.530 2258.435 2904.810 2258.805 ;
        RECT 13.890 2189.755 14.170 2190.125 ;
        RECT 13.960 2118.725 14.100 2189.755 ;
        RECT 13.890 2118.355 14.170 2118.725 ;
        RECT 13.960 1903.165 14.100 2118.355 ;
        RECT 2904.600 2082.685 2904.740 2258.435 ;
        RECT 2904.530 2082.315 2904.810 2082.685 ;
        RECT 2904.600 2024.205 2904.740 2082.315 ;
        RECT 2904.530 2023.835 2904.810 2024.205 ;
        RECT 13.890 1902.795 14.170 1903.165 ;
        RECT 13.960 1835.165 14.100 1902.795 ;
        RECT 2904.600 1848.085 2904.740 2023.835 ;
        RECT 2904.530 1847.715 2904.810 1848.085 ;
        RECT 13.890 1834.795 14.170 1835.165 ;
        RECT 17.110 1834.795 17.390 1835.165 ;
        RECT 17.180 1831.085 17.320 1834.795 ;
        RECT 17.110 1830.715 17.390 1831.085 ;
        RECT 17.180 1691.490 17.320 1830.715 ;
        RECT 2904.600 1789.605 2904.740 1847.715 ;
        RECT 2901.310 1789.235 2901.590 1789.605 ;
        RECT 2904.530 1789.235 2904.810 1789.605 ;
        RECT 17.120 1691.170 17.380 1691.490 ;
        RECT 17.180 1615.525 17.320 1691.170 ;
        RECT 2901.380 1690.810 2901.520 1789.235 ;
        RECT 2901.320 1690.490 2901.580 1690.810 ;
        RECT 13.890 1615.155 14.170 1615.525 ;
        RECT 17.110 1615.155 17.390 1615.525 ;
        RECT 13.960 1544.125 14.100 1615.155 ;
        RECT 2901.380 1613.485 2901.520 1690.490 ;
        RECT 2901.310 1613.115 2901.590 1613.485 ;
        RECT 2904.530 1613.115 2904.810 1613.485 ;
        RECT 2904.600 1554.325 2904.740 1613.115 ;
        RECT 2904.530 1553.955 2904.810 1554.325 ;
        RECT 13.890 1543.755 14.170 1544.125 ;
        RECT 13.960 1400.645 14.100 1543.755 ;
        RECT 13.890 1400.275 14.170 1400.645 ;
        RECT 13.960 1328.565 14.100 1400.275 ;
        RECT 2904.600 1378.885 2904.740 1553.955 ;
        RECT 2904.530 1378.515 2904.810 1378.885 ;
        RECT 13.890 1328.195 14.170 1328.565 ;
        RECT 13.960 1185.085 14.100 1328.195 ;
        RECT 2904.600 1319.725 2904.740 1378.515 ;
        RECT 2904.530 1319.355 2904.810 1319.725 ;
        RECT 13.890 1184.715 14.170 1185.085 ;
        RECT 13.960 1113.005 14.100 1184.715 ;
        RECT 2904.600 1144.285 2904.740 1319.355 ;
        RECT 2904.530 1143.915 2904.810 1144.285 ;
        RECT 13.890 1112.635 14.170 1113.005 ;
        RECT 13.960 969.525 14.100 1112.635 ;
        RECT 2904.600 1085.125 2904.740 1143.915 ;
        RECT 2904.530 1084.755 2904.810 1085.125 ;
        RECT 13.890 969.155 14.170 969.525 ;
        RECT 13.960 897.445 14.100 969.155 ;
        RECT 2904.600 909.685 2904.740 1084.755 ;
        RECT 2904.530 909.315 2904.810 909.685 ;
        RECT 13.890 897.075 14.170 897.445 ;
        RECT 13.960 753.965 14.100 897.075 ;
        RECT 2904.600 850.525 2904.740 909.315 ;
        RECT 2904.530 850.155 2904.810 850.525 ;
        RECT 13.890 753.595 14.170 753.965 ;
        RECT 13.960 681.885 14.100 753.595 ;
        RECT 13.890 681.515 14.170 681.885 ;
        RECT 13.960 538.405 14.100 681.515 ;
        RECT 2904.600 674.405 2904.740 850.155 ;
        RECT 2904.530 674.035 2904.810 674.405 ;
        RECT 2904.600 615.925 2904.740 674.035 ;
        RECT 2904.530 615.555 2904.810 615.925 ;
        RECT 13.890 538.035 14.170 538.405 ;
        RECT 13.960 466.325 14.100 538.035 ;
        RECT 13.890 465.955 14.170 466.325 ;
        RECT 13.960 322.845 14.100 465.955 ;
        RECT 2904.600 439.805 2904.740 615.555 ;
        RECT 2904.530 439.435 2904.810 439.805 ;
        RECT 2904.600 381.325 2904.740 439.435 ;
        RECT 2904.530 380.955 2904.810 381.325 ;
        RECT 13.890 322.475 14.170 322.845 ;
        RECT 13.960 250.765 14.100 322.475 ;
        RECT 13.890 250.395 14.170 250.765 ;
        RECT 13.960 107.285 14.100 250.395 ;
        RECT 2904.600 205.205 2904.740 380.955 ;
        RECT 2904.530 204.835 2904.810 205.205 ;
        RECT 2904.600 146.725 2904.740 204.835 ;
        RECT 2904.530 146.355 2904.810 146.725 ;
        RECT 13.890 106.915 14.170 107.285 ;
        RECT 13.960 35.885 14.100 106.915 ;
        RECT 13.890 35.515 14.170 35.885 ;
      LAYER via2 ;
        RECT 2904.530 2551.560 2904.810 2551.840 ;
        RECT 2904.530 2493.080 2904.810 2493.360 ;
        RECT 13.890 2477.440 14.170 2477.720 ;
        RECT 13.890 2405.360 14.170 2405.640 ;
        RECT 2904.530 2316.960 2904.810 2317.240 ;
        RECT 2904.530 2258.480 2904.810 2258.760 ;
        RECT 13.890 2189.800 14.170 2190.080 ;
        RECT 13.890 2118.400 14.170 2118.680 ;
        RECT 2904.530 2082.360 2904.810 2082.640 ;
        RECT 2904.530 2023.880 2904.810 2024.160 ;
        RECT 13.890 1902.840 14.170 1903.120 ;
        RECT 2904.530 1847.760 2904.810 1848.040 ;
        RECT 13.890 1834.840 14.170 1835.120 ;
        RECT 17.110 1834.840 17.390 1835.120 ;
        RECT 17.110 1830.760 17.390 1831.040 ;
        RECT 2901.310 1789.280 2901.590 1789.560 ;
        RECT 2904.530 1789.280 2904.810 1789.560 ;
        RECT 13.890 1615.200 14.170 1615.480 ;
        RECT 17.110 1615.200 17.390 1615.480 ;
        RECT 2901.310 1613.160 2901.590 1613.440 ;
        RECT 2904.530 1613.160 2904.810 1613.440 ;
        RECT 2904.530 1554.000 2904.810 1554.280 ;
        RECT 13.890 1543.800 14.170 1544.080 ;
        RECT 13.890 1400.320 14.170 1400.600 ;
        RECT 2904.530 1378.560 2904.810 1378.840 ;
        RECT 13.890 1328.240 14.170 1328.520 ;
        RECT 2904.530 1319.400 2904.810 1319.680 ;
        RECT 13.890 1184.760 14.170 1185.040 ;
        RECT 2904.530 1143.960 2904.810 1144.240 ;
        RECT 13.890 1112.680 14.170 1112.960 ;
        RECT 2904.530 1084.800 2904.810 1085.080 ;
        RECT 13.890 969.200 14.170 969.480 ;
        RECT 2904.530 909.360 2904.810 909.640 ;
        RECT 13.890 897.120 14.170 897.400 ;
        RECT 2904.530 850.200 2904.810 850.480 ;
        RECT 13.890 753.640 14.170 753.920 ;
        RECT 13.890 681.560 14.170 681.840 ;
        RECT 2904.530 674.080 2904.810 674.360 ;
        RECT 2904.530 615.600 2904.810 615.880 ;
        RECT 13.890 538.080 14.170 538.360 ;
        RECT 13.890 466.000 14.170 466.280 ;
        RECT 2904.530 439.480 2904.810 439.760 ;
        RECT 2904.530 381.000 2904.810 381.280 ;
        RECT 13.890 322.520 14.170 322.800 ;
        RECT 13.890 250.440 14.170 250.720 ;
        RECT 2904.530 204.880 2904.810 205.160 ;
        RECT 2904.530 146.400 2904.810 146.680 ;
        RECT 13.890 106.960 14.170 107.240 ;
        RECT 13.890 35.560 14.170 35.840 ;
      LAYER met3 ;
        RECT 2904.505 2551.850 2904.835 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2904.505 2551.550 2924.800 2551.850 ;
        RECT 2904.505 2551.535 2904.835 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 2904.505 2493.370 2904.835 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2904.505 2493.070 2924.800 2493.370 ;
        RECT 2904.505 2493.055 2904.835 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 13.865 2477.730 14.195 2477.745 ;
        RECT -4.800 2477.430 14.195 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 13.865 2477.415 14.195 2477.430 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 13.865 2405.650 14.195 2405.665 ;
        RECT -4.800 2405.350 14.195 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 13.865 2405.335 14.195 2405.350 ;
        RECT 2904.505 2317.250 2904.835 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2904.505 2316.950 2924.800 2317.250 ;
        RECT 2904.505 2316.935 2904.835 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 2904.505 2258.770 2904.835 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2904.505 2258.470 2924.800 2258.770 ;
        RECT 2904.505 2258.455 2904.835 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 13.865 2190.090 14.195 2190.105 ;
        RECT -4.800 2189.790 14.195 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 13.865 2189.775 14.195 2189.790 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 13.865 2118.690 14.195 2118.705 ;
        RECT -4.800 2118.390 14.195 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 13.865 2118.375 14.195 2118.390 ;
        RECT 2904.505 2082.650 2904.835 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2904.505 2082.350 2924.800 2082.650 ;
        RECT 2904.505 2082.335 2904.835 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 2904.505 2024.170 2904.835 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2904.505 2023.870 2924.800 2024.170 ;
        RECT 2904.505 2023.855 2904.835 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 13.865 1903.130 14.195 1903.145 ;
        RECT -4.800 1902.830 14.195 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 13.865 1902.815 14.195 1902.830 ;
        RECT 2904.505 1848.050 2904.835 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2904.505 1847.750 2924.800 1848.050 ;
        RECT 2904.505 1847.735 2904.835 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 13.865 1835.130 14.195 1835.145 ;
        RECT 17.085 1835.130 17.415 1835.145 ;
        RECT 13.865 1834.830 17.415 1835.130 ;
        RECT 13.865 1834.815 14.195 1834.830 ;
        RECT 17.085 1834.815 17.415 1834.830 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 17.085 1831.050 17.415 1831.065 ;
        RECT -4.800 1830.750 17.415 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 17.085 1830.735 17.415 1830.750 ;
        RECT 2901.285 1789.570 2901.615 1789.585 ;
        RECT 2904.505 1789.570 2904.835 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2901.285 1789.270 2924.800 1789.570 ;
        RECT 2901.285 1789.255 2901.615 1789.270 ;
        RECT 2904.505 1789.255 2904.835 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 13.865 1615.490 14.195 1615.505 ;
        RECT 17.085 1615.490 17.415 1615.505 ;
        RECT -4.800 1615.190 17.415 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 13.865 1615.175 14.195 1615.190 ;
        RECT 17.085 1615.175 17.415 1615.190 ;
        RECT 2901.285 1613.450 2901.615 1613.465 ;
        RECT 2904.505 1613.450 2904.835 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2901.285 1613.150 2924.800 1613.450 ;
        RECT 2901.285 1613.135 2901.615 1613.150 ;
        RECT 2904.505 1613.135 2904.835 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
        RECT 2904.505 1554.290 2904.835 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2904.505 1553.990 2924.800 1554.290 ;
        RECT 2904.505 1553.975 2904.835 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 13.865 1544.090 14.195 1544.105 ;
        RECT -4.800 1543.790 14.195 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 13.865 1543.775 14.195 1543.790 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 13.865 1400.610 14.195 1400.625 ;
        RECT -4.800 1400.310 14.195 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 13.865 1400.295 14.195 1400.310 ;
        RECT 2904.505 1378.850 2904.835 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2904.505 1378.550 2924.800 1378.850 ;
        RECT 2904.505 1378.535 2904.835 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 13.865 1328.530 14.195 1328.545 ;
        RECT -4.800 1328.230 14.195 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 13.865 1328.215 14.195 1328.230 ;
        RECT 2904.505 1319.690 2904.835 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2904.505 1319.390 2924.800 1319.690 ;
        RECT 2904.505 1319.375 2904.835 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 13.865 1185.050 14.195 1185.065 ;
        RECT -4.800 1184.750 14.195 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 13.865 1184.735 14.195 1184.750 ;
        RECT 2904.505 1144.250 2904.835 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2904.505 1143.950 2924.800 1144.250 ;
        RECT 2904.505 1143.935 2904.835 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 13.865 1112.970 14.195 1112.985 ;
        RECT -4.800 1112.670 14.195 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 13.865 1112.655 14.195 1112.670 ;
        RECT 2904.505 1085.090 2904.835 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2904.505 1084.790 2924.800 1085.090 ;
        RECT 2904.505 1084.775 2904.835 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 13.865 969.490 14.195 969.505 ;
        RECT -4.800 969.190 14.195 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 13.865 969.175 14.195 969.190 ;
        RECT 2904.505 909.650 2904.835 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2904.505 909.350 2924.800 909.650 ;
        RECT 2904.505 909.335 2904.835 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 13.865 897.410 14.195 897.425 ;
        RECT -4.800 897.110 14.195 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 13.865 897.095 14.195 897.110 ;
        RECT 2904.505 850.490 2904.835 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2904.505 850.190 2924.800 850.490 ;
        RECT 2904.505 850.175 2904.835 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 13.865 753.930 14.195 753.945 ;
        RECT -4.800 753.630 14.195 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 13.865 753.615 14.195 753.630 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 13.865 681.850 14.195 681.865 ;
        RECT -4.800 681.550 14.195 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 13.865 681.535 14.195 681.550 ;
        RECT 2904.505 674.370 2904.835 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2904.505 674.070 2924.800 674.370 ;
        RECT 2904.505 674.055 2904.835 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
        RECT 2904.505 615.890 2904.835 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2904.505 615.590 2924.800 615.890 ;
        RECT 2904.505 615.575 2904.835 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 13.865 538.370 14.195 538.385 ;
        RECT -4.800 538.070 14.195 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 13.865 538.055 14.195 538.070 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 13.865 466.290 14.195 466.305 ;
        RECT -4.800 465.990 14.195 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 13.865 465.975 14.195 465.990 ;
        RECT 2904.505 439.770 2904.835 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2904.505 439.470 2924.800 439.770 ;
        RECT 2904.505 439.455 2904.835 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
        RECT 2904.505 381.290 2904.835 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2904.505 380.990 2924.800 381.290 ;
        RECT 2904.505 380.975 2904.835 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 13.865 322.810 14.195 322.825 ;
        RECT -4.800 322.510 14.195 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 13.865 322.495 14.195 322.510 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 13.865 250.730 14.195 250.745 ;
        RECT -4.800 250.430 14.195 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 13.865 250.415 14.195 250.430 ;
        RECT 2904.505 205.170 2904.835 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2904.505 204.870 2924.800 205.170 ;
        RECT 2904.505 204.855 2904.835 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
        RECT 2904.505 146.690 2904.835 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2904.505 146.390 2924.800 146.690 ;
        RECT 2904.505 146.375 2904.835 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 13.865 107.250 14.195 107.265 ;
        RECT -4.800 106.950 14.195 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 13.865 106.935 14.195 106.950 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 13.865 35.850 14.195 35.865 ;
        RECT -4.800 35.550 14.195 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 13.865 35.535 14.195 35.550 ;
    END
  END io_oeb[0]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 6.510 324.600 6.830 324.660 ;
        RECT 6.510 324.460 54.000 324.600 ;
        RECT 6.510 324.400 6.830 324.460 ;
        RECT 2.830 17.580 3.150 17.640 ;
        RECT 6.510 17.580 6.830 17.640 ;
        RECT 2.830 17.440 6.830 17.580 ;
        RECT 2.830 17.380 3.150 17.440 ;
        RECT 6.510 17.380 6.830 17.440 ;
      LAYER via ;
        RECT 6.540 324.400 6.800 324.660 ;
        RECT 2.860 17.380 3.120 17.640 ;
        RECT 6.540 17.380 6.800 17.640 ;
      LAYER met2 ;
        RECT 6.540 324.370 6.800 324.690 ;
        RECT 6.600 17.670 6.740 324.370 ;
        RECT 2.860 17.350 3.120 17.670 ;
        RECT 6.540 17.350 6.800 17.670 ;
        RECT 2.920 2.400 3.060 17.350 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 13.410 338.200 13.730 338.260 ;
        RECT 13.410 338.060 54.000 338.200 ;
        RECT 13.410 338.000 13.730 338.060 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 13.410 17.580 13.730 17.640 ;
        RECT 8.350 17.440 13.730 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 13.410 17.380 13.730 17.440 ;
      LAYER via ;
        RECT 13.440 338.000 13.700 338.260 ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 13.440 17.380 13.700 17.640 ;
      LAYER met2 ;
        RECT 13.440 337.970 13.700 338.290 ;
        RECT 13.500 17.670 13.640 337.970 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 13.440 17.350 13.700 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.850 352.140 20.170 352.200 ;
        RECT 19.850 352.000 54.000 352.140 ;
        RECT 19.850 351.940 20.170 352.000 ;
        RECT 14.330 17.580 14.650 17.640 ;
        RECT 19.850 17.580 20.170 17.640 ;
        RECT 14.330 17.440 20.170 17.580 ;
        RECT 14.330 17.380 14.650 17.440 ;
        RECT 19.850 17.380 20.170 17.440 ;
      LAYER via ;
        RECT 19.880 351.940 20.140 352.200 ;
        RECT 14.360 17.380 14.620 17.640 ;
        RECT 19.880 17.380 20.140 17.640 ;
      LAYER met2 ;
        RECT 19.880 351.910 20.140 352.230 ;
        RECT 19.940 17.670 20.080 351.910 ;
        RECT 14.360 17.350 14.620 17.670 ;
        RECT 19.880 17.350 20.140 17.670 ;
        RECT 14.420 2.400 14.560 17.350 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 41.010 400.420 41.330 400.480 ;
        RECT 41.010 400.280 54.000 400.420 ;
        RECT 41.010 400.220 41.330 400.280 ;
        RECT 38.250 17.580 38.570 17.640 ;
        RECT 41.010 17.580 41.330 17.640 ;
        RECT 38.250 17.440 41.330 17.580 ;
        RECT 38.250 17.380 38.570 17.440 ;
        RECT 41.010 17.380 41.330 17.440 ;
      LAYER via ;
        RECT 41.040 400.220 41.300 400.480 ;
        RECT 38.280 17.380 38.540 17.640 ;
        RECT 41.040 17.380 41.300 17.640 ;
      LAYER met2 ;
        RECT 41.040 400.190 41.300 400.510 ;
        RECT 41.100 17.670 41.240 400.190 ;
        RECT 38.280 17.350 38.540 17.670 ;
        RECT 41.040 17.350 41.300 17.670 ;
        RECT 38.340 2.400 38.480 17.350 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 241.200 17.410 241.340 54.000 ;
        RECT 240.740 17.270 241.340 17.410 ;
        RECT 240.740 2.400 240.880 17.270 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 17.580 258.450 17.640 ;
        RECT 261.810 17.580 262.130 17.640 ;
        RECT 258.130 17.440 262.130 17.580 ;
        RECT 258.130 17.380 258.450 17.440 ;
        RECT 261.810 17.380 262.130 17.440 ;
      LAYER via ;
        RECT 258.160 17.380 258.420 17.640 ;
        RECT 261.840 17.380 262.100 17.640 ;
      LAYER met2 ;
        RECT 261.900 17.670 262.040 54.000 ;
        RECT 258.160 17.350 258.420 17.670 ;
        RECT 261.840 17.350 262.100 17.670 ;
        RECT 258.220 2.400 258.360 17.350 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 276.070 17.920 276.390 17.980 ;
        RECT 282.050 17.920 282.370 17.980 ;
        RECT 276.070 17.780 282.370 17.920 ;
        RECT 276.070 17.720 276.390 17.780 ;
        RECT 282.050 17.720 282.370 17.780 ;
      LAYER via ;
        RECT 276.100 17.720 276.360 17.980 ;
        RECT 282.080 17.720 282.340 17.980 ;
      LAYER met2 ;
        RECT 282.140 18.010 282.280 54.000 ;
        RECT 276.100 17.690 276.360 18.010 ;
        RECT 282.080 17.690 282.340 18.010 ;
        RECT 276.160 2.400 276.300 17.690 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 17.580 294.330 17.640 ;
        RECT 296.310 17.580 296.630 17.640 ;
        RECT 294.010 17.440 296.630 17.580 ;
        RECT 294.010 17.380 294.330 17.440 ;
        RECT 296.310 17.380 296.630 17.440 ;
      LAYER via ;
        RECT 294.040 17.380 294.300 17.640 ;
        RECT 296.340 17.380 296.600 17.640 ;
      LAYER met2 ;
        RECT 296.400 17.670 296.540 54.000 ;
        RECT 294.040 17.350 294.300 17.670 ;
        RECT 296.340 17.350 296.600 17.670 ;
        RECT 294.100 2.400 294.240 17.350 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 17.580 312.270 17.640 ;
        RECT 317.010 17.580 317.330 17.640 ;
        RECT 311.950 17.440 317.330 17.580 ;
        RECT 311.950 17.380 312.270 17.440 ;
        RECT 317.010 17.380 317.330 17.440 ;
      LAYER via ;
        RECT 311.980 17.380 312.240 17.640 ;
        RECT 317.040 17.380 317.300 17.640 ;
      LAYER met2 ;
        RECT 317.100 17.670 317.240 54.000 ;
        RECT 311.980 17.350 312.240 17.670 ;
        RECT 317.040 17.350 317.300 17.670 ;
        RECT 312.040 2.400 312.180 17.350 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 330.900 17.410 331.040 54.000 ;
        RECT 329.980 17.270 331.040 17.410 ;
        RECT 329.980 2.400 330.120 17.270 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 17.580 347.690 17.640 ;
        RECT 351.510 17.580 351.830 17.640 ;
        RECT 347.370 17.440 351.830 17.580 ;
        RECT 347.370 17.380 347.690 17.440 ;
        RECT 351.510 17.380 351.830 17.440 ;
      LAYER via ;
        RECT 347.400 17.380 347.660 17.640 ;
        RECT 351.540 17.380 351.800 17.640 ;
      LAYER met2 ;
        RECT 351.600 17.670 351.740 54.000 ;
        RECT 347.400 17.350 347.660 17.670 ;
        RECT 351.540 17.350 351.800 17.670 ;
        RECT 347.460 2.400 347.600 17.350 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.400 2.400 365.540 54.000 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 17.580 383.570 17.640 ;
        RECT 386.010 17.580 386.330 17.640 ;
        RECT 383.250 17.440 386.330 17.580 ;
        RECT 383.250 17.380 383.570 17.440 ;
        RECT 386.010 17.380 386.330 17.440 ;
      LAYER via ;
        RECT 383.280 17.380 383.540 17.640 ;
        RECT 386.040 17.380 386.300 17.640 ;
      LAYER met2 ;
        RECT 386.100 17.670 386.240 54.000 ;
        RECT 383.280 17.350 383.540 17.670 ;
        RECT 386.040 17.350 386.300 17.670 ;
        RECT 383.340 2.400 383.480 17.350 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 17.580 401.510 17.640 ;
        RECT 406.710 17.580 407.030 17.640 ;
        RECT 401.190 17.440 407.030 17.580 ;
        RECT 401.190 17.380 401.510 17.440 ;
        RECT 406.710 17.380 407.030 17.440 ;
      LAYER via ;
        RECT 401.220 17.380 401.480 17.640 ;
        RECT 406.740 17.380 407.000 17.640 ;
      LAYER met2 ;
        RECT 406.800 17.670 406.940 54.000 ;
        RECT 401.220 17.350 401.480 17.670 ;
        RECT 406.740 17.350 407.000 17.670 ;
        RECT 401.280 2.400 401.420 17.350 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 62.170 17.920 62.490 17.980 ;
        RECT 68.150 17.920 68.470 17.980 ;
        RECT 62.170 17.780 68.470 17.920 ;
        RECT 62.170 17.720 62.490 17.780 ;
        RECT 68.150 17.720 68.470 17.780 ;
      LAYER via ;
        RECT 62.200 17.720 62.460 17.980 ;
        RECT 68.180 17.720 68.440 17.980 ;
      LAYER met2 ;
        RECT 68.240 18.010 68.380 54.000 ;
        RECT 62.200 17.690 62.460 18.010 ;
        RECT 68.180 17.690 68.440 18.010 ;
        RECT 62.260 2.400 62.400 17.690 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 420.600 17.410 420.740 54.000 ;
        RECT 419.220 17.270 420.740 17.410 ;
        RECT 419.220 2.400 419.360 17.270 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 17.580 436.930 17.640 ;
        RECT 441.210 17.580 441.530 17.640 ;
        RECT 436.610 17.440 441.530 17.580 ;
        RECT 436.610 17.380 436.930 17.440 ;
        RECT 441.210 17.380 441.530 17.440 ;
      LAYER via ;
        RECT 436.640 17.380 436.900 17.640 ;
        RECT 441.240 17.380 441.500 17.640 ;
      LAYER met2 ;
        RECT 441.300 17.670 441.440 54.000 ;
        RECT 436.640 17.350 436.900 17.670 ;
        RECT 441.240 17.350 441.500 17.670 ;
        RECT 436.700 2.400 436.840 17.350 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 455.100 17.410 455.240 54.000 ;
        RECT 454.640 17.270 455.240 17.410 ;
        RECT 454.640 2.400 454.780 17.270 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.490 17.580 472.810 17.640 ;
        RECT 475.710 17.580 476.030 17.640 ;
        RECT 472.490 17.440 476.030 17.580 ;
        RECT 472.490 17.380 472.810 17.440 ;
        RECT 475.710 17.380 476.030 17.440 ;
      LAYER via ;
        RECT 472.520 17.380 472.780 17.640 ;
        RECT 475.740 17.380 476.000 17.640 ;
      LAYER met2 ;
        RECT 475.800 17.670 475.940 54.000 ;
        RECT 472.520 17.350 472.780 17.670 ;
        RECT 475.740 17.350 476.000 17.670 ;
        RECT 472.580 2.400 472.720 17.350 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 490.430 15.200 490.750 15.260 ;
        RECT 495.950 15.200 496.270 15.260 ;
        RECT 490.430 15.060 496.270 15.200 ;
        RECT 490.430 15.000 490.750 15.060 ;
        RECT 495.950 15.000 496.270 15.060 ;
      LAYER via ;
        RECT 490.460 15.000 490.720 15.260 ;
        RECT 495.980 15.000 496.240 15.260 ;
      LAYER met2 ;
        RECT 496.040 15.290 496.180 54.000 ;
        RECT 490.460 14.970 490.720 15.290 ;
        RECT 495.980 14.970 496.240 15.290 ;
        RECT 490.520 2.400 490.660 14.970 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 17.580 508.230 17.640 ;
        RECT 510.210 17.580 510.530 17.640 ;
        RECT 507.910 17.440 510.530 17.580 ;
        RECT 507.910 17.380 508.230 17.440 ;
        RECT 510.210 17.380 510.530 17.440 ;
      LAYER via ;
        RECT 507.940 17.380 508.200 17.640 ;
        RECT 510.240 17.380 510.500 17.640 ;
      LAYER met2 ;
        RECT 510.300 17.670 510.440 54.000 ;
        RECT 507.940 17.350 508.200 17.670 ;
        RECT 510.240 17.350 510.500 17.670 ;
        RECT 508.000 2.400 508.140 17.350 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 525.850 17.580 526.170 17.640 ;
        RECT 530.910 17.580 531.230 17.640 ;
        RECT 525.850 17.440 531.230 17.580 ;
        RECT 525.850 17.380 526.170 17.440 ;
        RECT 530.910 17.380 531.230 17.440 ;
      LAYER via ;
        RECT 525.880 17.380 526.140 17.640 ;
        RECT 530.940 17.380 531.200 17.640 ;
      LAYER met2 ;
        RECT 531.000 17.670 531.140 54.000 ;
        RECT 525.880 17.350 526.140 17.670 ;
        RECT 530.940 17.350 531.200 17.670 ;
        RECT 525.940 2.400 526.080 17.350 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 544.800 17.410 544.940 54.000 ;
        RECT 543.880 17.270 544.940 17.410 ;
        RECT 543.880 2.400 544.020 17.270 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 17.580 562.050 17.640 ;
        RECT 565.410 17.580 565.730 17.640 ;
        RECT 561.730 17.440 565.730 17.580 ;
        RECT 561.730 17.380 562.050 17.440 ;
        RECT 565.410 17.380 565.730 17.440 ;
      LAYER via ;
        RECT 561.760 17.380 562.020 17.640 ;
        RECT 565.440 17.380 565.700 17.640 ;
      LAYER met2 ;
        RECT 565.500 17.670 565.640 54.000 ;
        RECT 561.760 17.350 562.020 17.670 ;
        RECT 565.440 17.350 565.700 17.670 ;
        RECT 561.820 2.400 561.960 17.350 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.670 17.920 579.990 17.980 ;
        RECT 585.650 17.920 585.970 17.980 ;
        RECT 579.670 17.780 585.970 17.920 ;
        RECT 579.670 17.720 579.990 17.780 ;
        RECT 585.650 17.720 585.970 17.780 ;
      LAYER via ;
        RECT 579.700 17.720 579.960 17.980 ;
        RECT 585.680 17.720 585.940 17.980 ;
      LAYER met2 ;
        RECT 585.740 18.010 585.880 54.000 ;
        RECT 579.700 17.690 579.960 18.010 ;
        RECT 585.680 17.690 585.940 18.010 ;
        RECT 579.760 2.400 579.900 17.690 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 17.580 86.410 17.640 ;
        RECT 89.310 17.580 89.630 17.640 ;
        RECT 86.090 17.440 89.630 17.580 ;
        RECT 86.090 17.380 86.410 17.440 ;
        RECT 89.310 17.380 89.630 17.440 ;
      LAYER via ;
        RECT 86.120 17.380 86.380 17.640 ;
        RECT 89.340 17.380 89.600 17.640 ;
      LAYER met2 ;
        RECT 89.400 17.670 89.540 54.000 ;
        RECT 86.120 17.350 86.380 17.670 ;
        RECT 89.340 17.350 89.600 17.670 ;
        RECT 86.180 2.400 86.320 17.350 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 597.150 17.580 597.470 17.640 ;
        RECT 599.910 17.580 600.230 17.640 ;
        RECT 597.150 17.440 600.230 17.580 ;
        RECT 597.150 17.380 597.470 17.440 ;
        RECT 599.910 17.380 600.230 17.440 ;
      LAYER via ;
        RECT 597.180 17.380 597.440 17.640 ;
        RECT 599.940 17.380 600.200 17.640 ;
      LAYER met2 ;
        RECT 600.000 17.670 600.140 54.000 ;
        RECT 597.180 17.350 597.440 17.670 ;
        RECT 599.940 17.350 600.200 17.670 ;
        RECT 597.240 2.400 597.380 17.350 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 615.090 16.220 615.410 16.280 ;
        RECT 620.610 16.220 620.930 16.280 ;
        RECT 615.090 16.080 620.930 16.220 ;
        RECT 615.090 16.020 615.410 16.080 ;
        RECT 620.610 16.020 620.930 16.080 ;
      LAYER via ;
        RECT 615.120 16.020 615.380 16.280 ;
        RECT 620.640 16.020 620.900 16.280 ;
      LAYER met2 ;
        RECT 620.700 16.310 620.840 54.000 ;
        RECT 615.120 15.990 615.380 16.310 ;
        RECT 620.640 15.990 620.900 16.310 ;
        RECT 615.180 2.400 615.320 15.990 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.100 17.410 110.240 54.000 ;
        RECT 109.640 17.270 110.240 17.410 ;
        RECT 109.640 2.400 109.780 17.270 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 133.470 17.580 133.790 17.640 ;
        RECT 137.610 17.580 137.930 17.640 ;
        RECT 133.470 17.440 137.930 17.580 ;
        RECT 133.470 17.380 133.790 17.440 ;
        RECT 137.610 17.380 137.930 17.440 ;
      LAYER via ;
        RECT 133.500 17.380 133.760 17.640 ;
        RECT 137.640 17.380 137.900 17.640 ;
      LAYER met2 ;
        RECT 137.700 17.670 137.840 54.000 ;
        RECT 133.500 17.350 133.760 17.670 ;
        RECT 137.640 17.350 137.900 17.670 ;
        RECT 133.560 2.400 133.700 17.350 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.500 2.400 151.640 54.000 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 169.350 17.580 169.670 17.640 ;
        RECT 172.110 17.580 172.430 17.640 ;
        RECT 169.350 17.440 172.430 17.580 ;
        RECT 169.350 17.380 169.670 17.440 ;
        RECT 172.110 17.380 172.430 17.440 ;
      LAYER via ;
        RECT 169.380 17.380 169.640 17.640 ;
        RECT 172.140 17.380 172.400 17.640 ;
      LAYER met2 ;
        RECT 172.200 17.670 172.340 54.000 ;
        RECT 169.380 17.350 169.640 17.670 ;
        RECT 172.140 17.350 172.400 17.670 ;
        RECT 169.440 2.400 169.580 17.350 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 17.580 187.150 17.640 ;
        RECT 192.350 17.580 192.670 17.640 ;
        RECT 186.830 17.440 192.670 17.580 ;
        RECT 186.830 17.380 187.150 17.440 ;
        RECT 192.350 17.380 192.670 17.440 ;
      LAYER via ;
        RECT 186.860 17.380 187.120 17.640 ;
        RECT 192.380 17.380 192.640 17.640 ;
      LAYER met2 ;
        RECT 192.440 17.670 192.580 54.000 ;
        RECT 186.860 17.350 187.120 17.670 ;
        RECT 192.380 17.350 192.640 17.670 ;
        RECT 186.920 2.400 187.060 17.350 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.700 17.410 206.840 54.000 ;
        RECT 204.860 17.270 206.840 17.410 ;
        RECT 204.860 2.400 205.000 17.270 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 222.710 17.580 223.030 17.640 ;
        RECT 227.310 17.580 227.630 17.640 ;
        RECT 222.710 17.440 227.630 17.580 ;
        RECT 222.710 17.380 223.030 17.440 ;
        RECT 227.310 17.380 227.630 17.440 ;
      LAYER via ;
        RECT 222.740 17.380 223.000 17.640 ;
        RECT 227.340 17.380 227.600 17.640 ;
      LAYER met2 ;
        RECT 227.400 17.670 227.540 54.000 ;
        RECT 222.740 17.350 223.000 17.670 ;
        RECT 227.340 17.350 227.600 17.670 ;
        RECT 222.800 2.400 222.940 17.350 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 358.940 20.630 359.000 ;
        RECT 20.310 358.800 54.000 358.940 ;
        RECT 20.310 358.740 20.630 358.800 ;
      LAYER via ;
        RECT 20.340 358.740 20.600 359.000 ;
      LAYER met2 ;
        RECT 20.340 358.710 20.600 359.030 ;
        RECT 20.400 2.400 20.540 358.710 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.910 414.360 48.230 414.420 ;
        RECT 47.910 414.220 54.000 414.360 ;
        RECT 47.910 414.160 48.230 414.220 ;
        RECT 44.230 17.580 44.550 17.640 ;
        RECT 47.910 17.580 48.230 17.640 ;
        RECT 44.230 17.440 48.230 17.580 ;
        RECT 44.230 17.380 44.550 17.440 ;
        RECT 47.910 17.380 48.230 17.440 ;
      LAYER via ;
        RECT 47.940 414.160 48.200 414.420 ;
        RECT 44.260 17.380 44.520 17.640 ;
        RECT 47.940 17.380 48.200 17.640 ;
      LAYER met2 ;
        RECT 47.940 414.130 48.200 414.450 ;
        RECT 48.000 17.670 48.140 414.130 ;
        RECT 44.260 17.350 44.520 17.670 ;
        RECT 47.940 17.350 48.200 17.670 ;
        RECT 44.320 2.400 44.460 17.350 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 248.100 17.580 248.240 54.000 ;
        RECT 246.720 17.440 248.240 17.580 ;
        RECT 246.720 2.400 246.860 17.440 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 264.110 15.200 264.430 15.260 ;
        RECT 268.710 15.200 269.030 15.260 ;
        RECT 264.110 15.060 269.030 15.200 ;
        RECT 264.110 15.000 264.430 15.060 ;
        RECT 268.710 15.000 269.030 15.060 ;
      LAYER via ;
        RECT 264.140 15.000 264.400 15.260 ;
        RECT 268.740 15.000 269.000 15.260 ;
      LAYER met2 ;
        RECT 268.800 15.290 268.940 54.000 ;
        RECT 264.140 14.970 264.400 15.290 ;
        RECT 268.740 14.970 269.000 15.290 ;
        RECT 264.200 2.400 264.340 14.970 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.600 17.410 282.740 54.000 ;
        RECT 282.140 17.270 282.740 17.410 ;
        RECT 282.140 2.400 282.280 17.270 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 299.990 15.200 300.310 15.260 ;
        RECT 303.210 15.200 303.530 15.260 ;
        RECT 299.990 15.060 303.530 15.200 ;
        RECT 299.990 15.000 300.310 15.060 ;
        RECT 303.210 15.000 303.530 15.060 ;
      LAYER via ;
        RECT 300.020 15.000 300.280 15.260 ;
        RECT 303.240 15.000 303.500 15.260 ;
      LAYER met2 ;
        RECT 303.300 15.290 303.440 54.000 ;
        RECT 300.020 14.970 300.280 15.290 ;
        RECT 303.240 14.970 303.500 15.290 ;
        RECT 300.080 2.400 300.220 14.970 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.930 17.580 318.250 17.640 ;
        RECT 323.450 17.580 323.770 17.640 ;
        RECT 317.930 17.440 323.770 17.580 ;
        RECT 317.930 17.380 318.250 17.440 ;
        RECT 323.450 17.380 323.770 17.440 ;
      LAYER via ;
        RECT 317.960 17.380 318.220 17.640 ;
        RECT 323.480 17.380 323.740 17.640 ;
      LAYER met2 ;
        RECT 323.540 17.670 323.680 54.000 ;
        RECT 317.960 17.350 318.220 17.670 ;
        RECT 323.480 17.350 323.740 17.670 ;
        RECT 318.020 2.400 318.160 17.350 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 337.800 17.410 337.940 54.000 ;
        RECT 335.960 17.270 337.940 17.410 ;
        RECT 335.960 2.400 336.100 17.270 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 353.350 17.580 353.670 17.640 ;
        RECT 358.410 17.580 358.730 17.640 ;
        RECT 353.350 17.440 358.730 17.580 ;
        RECT 353.350 17.380 353.670 17.440 ;
        RECT 358.410 17.380 358.730 17.440 ;
      LAYER via ;
        RECT 353.380 17.380 353.640 17.640 ;
        RECT 358.440 17.380 358.700 17.640 ;
      LAYER met2 ;
        RECT 358.500 17.670 358.640 54.000 ;
        RECT 353.380 17.350 353.640 17.670 ;
        RECT 358.440 17.350 358.700 17.670 ;
        RECT 353.440 2.400 353.580 17.350 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 372.300 17.410 372.440 54.000 ;
        RECT 371.380 17.270 372.440 17.410 ;
        RECT 371.380 2.400 371.520 17.270 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 389.230 17.580 389.550 17.640 ;
        RECT 392.910 17.580 393.230 17.640 ;
        RECT 389.230 17.440 393.230 17.580 ;
        RECT 389.230 17.380 389.550 17.440 ;
        RECT 392.910 17.380 393.230 17.440 ;
      LAYER via ;
        RECT 389.260 17.380 389.520 17.640 ;
        RECT 392.940 17.380 393.200 17.640 ;
      LAYER met2 ;
        RECT 393.000 17.670 393.140 54.000 ;
        RECT 389.260 17.350 389.520 17.670 ;
        RECT 392.940 17.350 393.200 17.670 ;
        RECT 389.320 2.400 389.460 17.350 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 407.170 17.920 407.490 17.980 ;
        RECT 413.150 17.920 413.470 17.980 ;
        RECT 407.170 17.780 413.470 17.920 ;
        RECT 407.170 17.720 407.490 17.780 ;
        RECT 413.150 17.720 413.470 17.780 ;
      LAYER via ;
        RECT 407.200 17.720 407.460 17.980 ;
        RECT 413.180 17.720 413.440 17.980 ;
      LAYER met2 ;
        RECT 413.240 18.010 413.380 54.000 ;
        RECT 407.200 17.690 407.460 18.010 ;
        RECT 413.180 17.690 413.440 18.010 ;
        RECT 407.260 2.400 407.400 17.690 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.700 17.410 68.840 54.000 ;
        RECT 68.240 17.270 68.840 17.410 ;
        RECT 68.240 2.400 68.380 17.270 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 424.650 17.580 424.970 17.640 ;
        RECT 427.410 17.580 427.730 17.640 ;
        RECT 424.650 17.440 427.730 17.580 ;
        RECT 424.650 17.380 424.970 17.440 ;
        RECT 427.410 17.380 427.730 17.440 ;
      LAYER via ;
        RECT 424.680 17.380 424.940 17.640 ;
        RECT 427.440 17.380 427.700 17.640 ;
      LAYER met2 ;
        RECT 427.500 17.670 427.640 54.000 ;
        RECT 424.680 17.350 424.940 17.670 ;
        RECT 427.440 17.350 427.700 17.670 ;
        RECT 424.740 2.400 424.880 17.350 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 442.590 17.580 442.910 17.640 ;
        RECT 448.110 17.580 448.430 17.640 ;
        RECT 442.590 17.440 448.430 17.580 ;
        RECT 442.590 17.380 442.910 17.440 ;
        RECT 448.110 17.380 448.430 17.440 ;
      LAYER via ;
        RECT 442.620 17.380 442.880 17.640 ;
        RECT 448.140 17.380 448.400 17.640 ;
      LAYER met2 ;
        RECT 448.200 17.670 448.340 54.000 ;
        RECT 442.620 17.350 442.880 17.670 ;
        RECT 448.140 17.350 448.400 17.670 ;
        RECT 442.680 2.400 442.820 17.350 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 462.000 17.410 462.140 54.000 ;
        RECT 460.620 17.270 462.140 17.410 ;
        RECT 460.620 2.400 460.760 17.270 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 478.470 17.580 478.790 17.640 ;
        RECT 482.610 17.580 482.930 17.640 ;
        RECT 478.470 17.440 482.930 17.580 ;
        RECT 478.470 17.380 478.790 17.440 ;
        RECT 482.610 17.380 482.930 17.440 ;
      LAYER via ;
        RECT 478.500 17.380 478.760 17.640 ;
        RECT 482.640 17.380 482.900 17.640 ;
      LAYER met2 ;
        RECT 482.700 17.670 482.840 54.000 ;
        RECT 478.500 17.350 478.760 17.670 ;
        RECT 482.640 17.350 482.900 17.670 ;
        RECT 478.560 2.400 478.700 17.350 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.500 2.400 496.640 54.000 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 513.890 17.580 514.210 17.640 ;
        RECT 517.110 17.580 517.430 17.640 ;
        RECT 513.890 17.440 517.430 17.580 ;
        RECT 513.890 17.380 514.210 17.440 ;
        RECT 517.110 17.380 517.430 17.440 ;
      LAYER via ;
        RECT 513.920 17.380 514.180 17.640 ;
        RECT 517.140 17.380 517.400 17.640 ;
      LAYER met2 ;
        RECT 517.200 17.670 517.340 54.000 ;
        RECT 513.920 17.350 514.180 17.670 ;
        RECT 517.140 17.350 517.400 17.670 ;
        RECT 513.980 2.400 514.120 17.350 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 531.830 15.200 532.150 15.260 ;
        RECT 537.350 15.200 537.670 15.260 ;
        RECT 531.830 15.060 537.670 15.200 ;
        RECT 531.830 15.000 532.150 15.060 ;
        RECT 537.350 15.000 537.670 15.060 ;
      LAYER via ;
        RECT 531.860 15.000 532.120 15.260 ;
        RECT 537.380 15.000 537.640 15.260 ;
      LAYER met2 ;
        RECT 537.440 15.290 537.580 54.000 ;
        RECT 531.860 14.970 532.120 15.290 ;
        RECT 537.380 14.970 537.640 15.290 ;
        RECT 531.920 2.400 532.060 14.970 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 551.700 17.410 551.840 54.000 ;
        RECT 549.860 17.270 551.840 17.410 ;
        RECT 549.860 2.400 550.000 17.270 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 567.710 17.580 568.030 17.640 ;
        RECT 572.310 17.580 572.630 17.640 ;
        RECT 567.710 17.440 572.630 17.580 ;
        RECT 567.710 17.380 568.030 17.440 ;
        RECT 572.310 17.380 572.630 17.440 ;
      LAYER via ;
        RECT 567.740 17.380 568.000 17.640 ;
        RECT 572.340 17.380 572.600 17.640 ;
      LAYER met2 ;
        RECT 572.400 17.670 572.540 54.000 ;
        RECT 567.740 17.350 568.000 17.670 ;
        RECT 572.340 17.350 572.600 17.670 ;
        RECT 567.800 2.400 567.940 17.350 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 586.200 17.410 586.340 54.000 ;
        RECT 585.740 17.270 586.340 17.410 ;
        RECT 585.740 2.400 585.880 17.270 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 91.610 17.580 91.930 17.640 ;
        RECT 96.210 17.580 96.530 17.640 ;
        RECT 91.610 17.440 96.530 17.580 ;
        RECT 91.610 17.380 91.930 17.440 ;
        RECT 96.210 17.380 96.530 17.440 ;
      LAYER via ;
        RECT 91.640 17.380 91.900 17.640 ;
        RECT 96.240 17.380 96.500 17.640 ;
      LAYER met2 ;
        RECT 96.300 17.670 96.440 54.000 ;
        RECT 91.640 17.350 91.900 17.670 ;
        RECT 96.240 17.350 96.500 17.670 ;
        RECT 91.700 2.400 91.840 17.350 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 603.130 17.580 603.450 17.640 ;
        RECT 606.810 17.580 607.130 17.640 ;
        RECT 603.130 17.440 607.130 17.580 ;
        RECT 603.130 17.380 603.450 17.440 ;
        RECT 606.810 17.380 607.130 17.440 ;
      LAYER via ;
        RECT 603.160 17.380 603.420 17.640 ;
        RECT 606.840 17.380 607.100 17.640 ;
      LAYER met2 ;
        RECT 606.900 17.670 607.040 54.000 ;
        RECT 603.160 17.350 603.420 17.670 ;
        RECT 606.840 17.350 607.100 17.670 ;
        RECT 603.220 2.400 603.360 17.350 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 621.070 17.580 621.390 17.640 ;
        RECT 631.190 17.580 631.510 17.640 ;
        RECT 621.070 17.440 631.510 17.580 ;
        RECT 621.070 17.380 621.390 17.440 ;
        RECT 631.190 17.380 631.510 17.440 ;
      LAYER via ;
        RECT 621.100 17.380 621.360 17.640 ;
        RECT 631.220 17.380 631.480 17.640 ;
      LAYER met2 ;
        RECT 631.280 17.670 631.420 54.000 ;
        RECT 621.100 17.350 621.360 17.670 ;
        RECT 631.220 17.350 631.480 17.670 ;
        RECT 621.160 2.400 621.300 17.350 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.000 17.410 117.140 54.000 ;
        RECT 115.620 17.270 117.140 17.410 ;
        RECT 115.620 2.400 115.760 17.270 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 139.450 17.580 139.770 17.640 ;
        RECT 144.510 17.580 144.830 17.640 ;
        RECT 139.450 17.440 144.830 17.580 ;
        RECT 139.450 17.380 139.770 17.440 ;
        RECT 144.510 17.380 144.830 17.440 ;
      LAYER via ;
        RECT 139.480 17.380 139.740 17.640 ;
        RECT 144.540 17.380 144.800 17.640 ;
      LAYER met2 ;
        RECT 144.600 17.670 144.740 54.000 ;
        RECT 139.480 17.350 139.740 17.670 ;
        RECT 144.540 17.350 144.800 17.670 ;
        RECT 139.540 2.400 139.680 17.350 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 158.400 17.410 158.540 54.000 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 174.870 17.580 175.190 17.640 ;
        RECT 179.010 17.580 179.330 17.640 ;
        RECT 174.870 17.440 179.330 17.580 ;
        RECT 174.870 17.380 175.190 17.440 ;
        RECT 179.010 17.380 179.330 17.440 ;
      LAYER via ;
        RECT 174.900 17.380 175.160 17.640 ;
        RECT 179.040 17.380 179.300 17.640 ;
      LAYER met2 ;
        RECT 179.100 17.670 179.240 54.000 ;
        RECT 174.900 17.350 175.160 17.670 ;
        RECT 179.040 17.350 179.300 17.670 ;
        RECT 174.960 2.400 175.100 17.350 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.900 2.400 193.040 54.000 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 210.750 17.580 211.070 17.640 ;
        RECT 213.510 17.580 213.830 17.640 ;
        RECT 210.750 17.440 213.830 17.580 ;
        RECT 210.750 17.380 211.070 17.440 ;
        RECT 213.510 17.380 213.830 17.440 ;
      LAYER via ;
        RECT 210.780 17.380 211.040 17.640 ;
        RECT 213.540 17.380 213.800 17.640 ;
      LAYER met2 ;
        RECT 213.600 17.670 213.740 54.000 ;
        RECT 210.780 17.350 211.040 17.670 ;
        RECT 213.540 17.350 213.800 17.670 ;
        RECT 210.840 2.400 210.980 17.350 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 228.690 17.580 229.010 17.640 ;
        RECT 234.210 17.580 234.530 17.640 ;
        RECT 228.690 17.440 234.530 17.580 ;
        RECT 228.690 17.380 229.010 17.440 ;
        RECT 234.210 17.380 234.530 17.440 ;
      LAYER via ;
        RECT 228.720 17.380 228.980 17.640 ;
        RECT 234.240 17.380 234.500 17.640 ;
      LAYER met2 ;
        RECT 234.300 17.670 234.440 54.000 ;
        RECT 228.720 17.350 228.980 17.670 ;
        RECT 234.240 17.350 234.500 17.670 ;
        RECT 228.780 2.400 228.920 17.350 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 50.210 17.580 50.530 17.640 ;
        RECT 54.810 17.580 55.130 17.640 ;
        RECT 50.210 17.440 55.130 17.580 ;
        RECT 50.210 17.380 50.530 17.440 ;
        RECT 54.810 17.380 55.130 17.440 ;
      LAYER via ;
        RECT 50.240 17.380 50.500 17.640 ;
        RECT 54.840 17.380 55.100 17.640 ;
      LAYER met2 ;
        RECT 54.900 17.670 55.040 54.000 ;
        RECT 50.240 17.350 50.500 17.670 ;
        RECT 54.840 17.350 55.100 17.670 ;
        RECT 50.300 2.400 50.440 17.350 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 252.610 17.580 252.930 17.640 ;
        RECT 254.910 17.580 255.230 17.640 ;
        RECT 252.610 17.440 255.230 17.580 ;
        RECT 252.610 17.380 252.930 17.440 ;
        RECT 254.910 17.380 255.230 17.440 ;
      LAYER via ;
        RECT 252.640 17.380 252.900 17.640 ;
        RECT 254.940 17.380 255.200 17.640 ;
      LAYER met2 ;
        RECT 255.000 17.670 255.140 54.000 ;
        RECT 252.640 17.350 252.900 17.670 ;
        RECT 254.940 17.350 255.200 17.670 ;
        RECT 252.700 2.400 252.840 17.350 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 270.090 17.580 270.410 17.640 ;
        RECT 275.610 17.580 275.930 17.640 ;
        RECT 270.090 17.440 275.930 17.580 ;
        RECT 270.090 17.380 270.410 17.440 ;
        RECT 275.610 17.380 275.930 17.440 ;
      LAYER via ;
        RECT 270.120 17.380 270.380 17.640 ;
        RECT 275.640 17.380 275.900 17.640 ;
      LAYER met2 ;
        RECT 275.700 17.670 275.840 54.000 ;
        RECT 270.120 17.350 270.380 17.670 ;
        RECT 275.640 17.350 275.900 17.670 ;
        RECT 270.180 2.400 270.320 17.350 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 289.500 17.410 289.640 54.000 ;
        RECT 288.120 17.270 289.640 17.410 ;
        RECT 288.120 2.400 288.260 17.270 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 305.970 17.580 306.290 17.640 ;
        RECT 310.110 17.580 310.430 17.640 ;
        RECT 305.970 17.440 310.430 17.580 ;
        RECT 305.970 17.380 306.290 17.440 ;
        RECT 310.110 17.380 310.430 17.440 ;
      LAYER via ;
        RECT 306.000 17.380 306.260 17.640 ;
        RECT 310.140 17.380 310.400 17.640 ;
      LAYER met2 ;
        RECT 310.200 17.670 310.340 54.000 ;
        RECT 306.000 17.350 306.260 17.670 ;
        RECT 310.140 17.350 310.400 17.670 ;
        RECT 306.060 2.400 306.200 17.350 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 324.000 2.400 324.140 54.000 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 341.390 15.200 341.710 15.260 ;
        RECT 344.610 15.200 344.930 15.260 ;
        RECT 341.390 15.060 344.930 15.200 ;
        RECT 341.390 15.000 341.710 15.060 ;
        RECT 344.610 15.000 344.930 15.060 ;
      LAYER via ;
        RECT 341.420 15.000 341.680 15.260 ;
        RECT 344.640 15.000 344.900 15.260 ;
      LAYER met2 ;
        RECT 344.700 15.290 344.840 54.000 ;
        RECT 341.420 14.970 341.680 15.290 ;
        RECT 344.640 14.970 344.900 15.290 ;
        RECT 341.480 2.400 341.620 14.970 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 359.330 17.580 359.650 17.640 ;
        RECT 364.850 17.580 365.170 17.640 ;
        RECT 359.330 17.440 365.170 17.580 ;
        RECT 359.330 17.380 359.650 17.440 ;
        RECT 364.850 17.380 365.170 17.440 ;
      LAYER via ;
        RECT 359.360 17.380 359.620 17.640 ;
        RECT 364.880 17.380 365.140 17.640 ;
      LAYER met2 ;
        RECT 364.940 17.670 365.080 54.000 ;
        RECT 359.360 17.350 359.620 17.670 ;
        RECT 364.880 17.350 365.140 17.670 ;
        RECT 359.420 2.400 359.560 17.350 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 379.200 17.410 379.340 54.000 ;
        RECT 377.360 17.270 379.340 17.410 ;
        RECT 377.360 2.400 377.500 17.270 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 395.210 17.580 395.530 17.640 ;
        RECT 399.810 17.580 400.130 17.640 ;
        RECT 395.210 17.440 400.130 17.580 ;
        RECT 395.210 17.380 395.530 17.440 ;
        RECT 399.810 17.380 400.130 17.440 ;
      LAYER via ;
        RECT 395.240 17.380 395.500 17.640 ;
        RECT 399.840 17.380 400.100 17.640 ;
      LAYER met2 ;
        RECT 399.900 17.670 400.040 54.000 ;
        RECT 395.240 17.350 395.500 17.670 ;
        RECT 399.840 17.350 400.100 17.670 ;
        RECT 395.300 2.400 395.440 17.350 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.700 17.410 413.840 54.000 ;
        RECT 413.240 17.270 413.840 17.410 ;
        RECT 413.240 2.400 413.380 17.270 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.600 17.410 75.740 54.000 ;
        RECT 74.220 17.270 75.740 17.410 ;
        RECT 74.220 2.400 74.360 17.270 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 430.630 17.580 430.950 17.640 ;
        RECT 434.310 17.580 434.630 17.640 ;
        RECT 430.630 17.440 434.630 17.580 ;
        RECT 430.630 17.380 430.950 17.440 ;
        RECT 434.310 17.380 434.630 17.440 ;
      LAYER via ;
        RECT 430.660 17.380 430.920 17.640 ;
        RECT 434.340 17.380 434.600 17.640 ;
      LAYER met2 ;
        RECT 434.400 17.670 434.540 54.000 ;
        RECT 430.660 17.350 430.920 17.670 ;
        RECT 434.340 17.350 434.600 17.670 ;
        RECT 430.720 2.400 430.860 17.350 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 448.570 17.920 448.890 17.980 ;
        RECT 454.550 17.920 454.870 17.980 ;
        RECT 448.570 17.780 454.870 17.920 ;
        RECT 448.570 17.720 448.890 17.780 ;
        RECT 454.550 17.720 454.870 17.780 ;
      LAYER via ;
        RECT 448.600 17.720 448.860 17.980 ;
        RECT 454.580 17.720 454.840 17.980 ;
      LAYER met2 ;
        RECT 454.640 18.010 454.780 54.000 ;
        RECT 448.600 17.690 448.860 18.010 ;
        RECT 454.580 17.690 454.840 18.010 ;
        RECT 448.660 2.400 448.800 17.690 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 466.510 16.900 466.830 16.960 ;
        RECT 468.810 16.900 469.130 16.960 ;
        RECT 466.510 16.760 469.130 16.900 ;
        RECT 466.510 16.700 466.830 16.760 ;
        RECT 468.810 16.700 469.130 16.760 ;
      LAYER via ;
        RECT 466.540 16.700 466.800 16.960 ;
        RECT 468.840 16.700 469.100 16.960 ;
      LAYER met2 ;
        RECT 468.900 16.990 469.040 54.000 ;
        RECT 466.540 16.670 466.800 16.990 ;
        RECT 468.840 16.670 469.100 16.990 ;
        RECT 466.600 2.400 466.740 16.670 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 484.450 16.560 484.770 16.620 ;
        RECT 489.510 16.560 489.830 16.620 ;
        RECT 484.450 16.420 489.830 16.560 ;
        RECT 484.450 16.360 484.770 16.420 ;
        RECT 489.510 16.360 489.830 16.420 ;
      LAYER via ;
        RECT 484.480 16.360 484.740 16.620 ;
        RECT 489.540 16.360 489.800 16.620 ;
      LAYER met2 ;
        RECT 489.600 16.650 489.740 54.000 ;
        RECT 484.480 16.330 484.740 16.650 ;
        RECT 489.540 16.330 489.800 16.650 ;
        RECT 484.540 2.400 484.680 16.330 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 503.400 17.410 503.540 54.000 ;
        RECT 502.480 17.270 503.540 17.410 ;
        RECT 502.480 2.400 502.620 17.270 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 519.870 17.580 520.190 17.640 ;
        RECT 524.010 17.580 524.330 17.640 ;
        RECT 519.870 17.440 524.330 17.580 ;
        RECT 519.870 17.380 520.190 17.440 ;
        RECT 524.010 17.380 524.330 17.440 ;
      LAYER via ;
        RECT 519.900 17.380 520.160 17.640 ;
        RECT 524.040 17.380 524.300 17.640 ;
      LAYER met2 ;
        RECT 524.100 17.670 524.240 54.000 ;
        RECT 519.900 17.350 520.160 17.670 ;
        RECT 524.040 17.350 524.300 17.670 ;
        RECT 519.960 2.400 520.100 17.350 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.900 2.400 538.040 54.000 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 555.750 17.580 556.070 17.640 ;
        RECT 558.510 17.580 558.830 17.640 ;
        RECT 555.750 17.440 558.830 17.580 ;
        RECT 555.750 17.380 556.070 17.440 ;
        RECT 558.510 17.380 558.830 17.440 ;
      LAYER via ;
        RECT 555.780 17.380 556.040 17.640 ;
        RECT 558.540 17.380 558.800 17.640 ;
      LAYER met2 ;
        RECT 558.600 17.670 558.740 54.000 ;
        RECT 555.780 17.350 556.040 17.670 ;
        RECT 558.540 17.350 558.800 17.670 ;
        RECT 555.840 2.400 555.980 17.350 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 573.690 15.200 574.010 15.260 ;
        RECT 579.210 15.200 579.530 15.260 ;
        RECT 573.690 15.060 579.530 15.200 ;
        RECT 573.690 15.000 574.010 15.060 ;
        RECT 579.210 15.000 579.530 15.060 ;
      LAYER via ;
        RECT 573.720 15.000 573.980 15.260 ;
        RECT 579.240 15.000 579.500 15.260 ;
      LAYER met2 ;
        RECT 579.300 15.290 579.440 54.000 ;
        RECT 573.720 14.970 573.980 15.290 ;
        RECT 579.240 14.970 579.500 15.290 ;
        RECT 573.780 2.400 573.920 14.970 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 593.100 17.410 593.240 54.000 ;
        RECT 591.260 17.270 593.240 17.410 ;
        RECT 591.260 2.400 591.400 17.270 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 97.590 16.560 97.910 16.620 ;
        RECT 103.110 16.560 103.430 16.620 ;
        RECT 97.590 16.420 103.430 16.560 ;
        RECT 97.590 16.360 97.910 16.420 ;
        RECT 103.110 16.360 103.430 16.420 ;
      LAYER via ;
        RECT 97.620 16.360 97.880 16.620 ;
        RECT 103.140 16.360 103.400 16.620 ;
      LAYER met2 ;
        RECT 103.200 16.650 103.340 54.000 ;
        RECT 97.620 16.330 97.880 16.650 ;
        RECT 103.140 16.330 103.400 16.650 ;
        RECT 97.680 2.400 97.820 16.330 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 609.110 17.580 609.430 17.640 ;
        RECT 613.710 17.580 614.030 17.640 ;
        RECT 609.110 17.440 614.030 17.580 ;
        RECT 609.110 17.380 609.430 17.440 ;
        RECT 613.710 17.380 614.030 17.440 ;
      LAYER via ;
        RECT 609.140 17.380 609.400 17.640 ;
        RECT 613.740 17.380 614.000 17.640 ;
      LAYER met2 ;
        RECT 613.800 17.670 613.940 54.000 ;
        RECT 609.140 17.350 609.400 17.670 ;
        RECT 613.740 17.350 614.000 17.670 ;
        RECT 609.200 2.400 609.340 17.350 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 627.600 3.130 627.740 54.000 ;
        RECT 627.140 2.990 627.740 3.130 ;
        RECT 627.140 2.400 627.280 2.990 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 17.580 121.830 17.640 ;
        RECT 123.810 17.580 124.130 17.640 ;
        RECT 121.510 17.440 124.130 17.580 ;
        RECT 121.510 17.380 121.830 17.440 ;
        RECT 123.810 17.380 124.130 17.440 ;
      LAYER via ;
        RECT 121.540 17.380 121.800 17.640 ;
        RECT 123.840 17.380 124.100 17.640 ;
      LAYER met2 ;
        RECT 123.900 17.670 124.040 54.000 ;
        RECT 121.540 17.350 121.800 17.670 ;
        RECT 123.840 17.350 124.100 17.670 ;
        RECT 121.600 2.400 121.740 17.350 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 145.430 15.200 145.750 15.260 ;
        RECT 150.950 15.200 151.270 15.260 ;
        RECT 145.430 15.060 151.270 15.200 ;
        RECT 145.430 15.000 145.750 15.060 ;
        RECT 150.950 15.000 151.270 15.060 ;
      LAYER via ;
        RECT 145.460 15.000 145.720 15.260 ;
        RECT 150.980 15.000 151.240 15.260 ;
      LAYER met2 ;
        RECT 151.040 15.290 151.180 54.000 ;
        RECT 145.460 14.970 145.720 15.290 ;
        RECT 150.980 14.970 151.240 15.290 ;
        RECT 145.520 2.400 145.660 14.970 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 165.300 17.410 165.440 54.000 ;
        RECT 163.460 17.270 165.440 17.410 ;
        RECT 163.460 2.400 163.600 17.270 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 180.850 17.580 181.170 17.640 ;
        RECT 185.910 17.580 186.230 17.640 ;
        RECT 180.850 17.440 186.230 17.580 ;
        RECT 180.850 17.380 181.170 17.440 ;
        RECT 185.910 17.380 186.230 17.440 ;
      LAYER via ;
        RECT 180.880 17.380 181.140 17.640 ;
        RECT 185.940 17.380 186.200 17.640 ;
      LAYER met2 ;
        RECT 186.000 17.670 186.140 54.000 ;
        RECT 180.880 17.350 181.140 17.670 ;
        RECT 185.940 17.350 186.200 17.670 ;
        RECT 180.940 2.400 181.080 17.350 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 199.800 17.410 199.940 54.000 ;
        RECT 198.880 17.270 199.940 17.410 ;
        RECT 198.880 2.400 199.020 17.270 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 216.730 17.580 217.050 17.640 ;
        RECT 220.410 17.580 220.730 17.640 ;
        RECT 216.730 17.440 220.730 17.580 ;
        RECT 216.730 17.380 217.050 17.440 ;
        RECT 220.410 17.380 220.730 17.440 ;
      LAYER via ;
        RECT 216.760 17.380 217.020 17.640 ;
        RECT 220.440 17.380 220.700 17.640 ;
      LAYER met2 ;
        RECT 220.500 17.670 220.640 54.000 ;
        RECT 216.760 17.350 217.020 17.670 ;
        RECT 220.440 17.350 220.700 17.670 ;
        RECT 216.820 2.400 216.960 17.350 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 234.670 17.920 234.990 17.980 ;
        RECT 240.650 17.920 240.970 17.980 ;
        RECT 234.670 17.780 240.970 17.920 ;
        RECT 234.670 17.720 234.990 17.780 ;
        RECT 240.650 17.720 240.970 17.780 ;
      LAYER via ;
        RECT 234.700 17.720 234.960 17.980 ;
        RECT 240.680 17.720 240.940 17.980 ;
      LAYER met2 ;
        RECT 240.740 18.010 240.880 54.000 ;
        RECT 234.700 17.690 234.960 18.010 ;
        RECT 240.680 17.690 240.940 18.010 ;
        RECT 234.760 2.400 234.900 17.690 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 56.190 17.580 56.510 17.640 ;
        RECT 61.710 17.580 62.030 17.640 ;
        RECT 56.190 17.440 62.030 17.580 ;
        RECT 56.190 17.380 56.510 17.440 ;
        RECT 61.710 17.380 62.030 17.440 ;
      LAYER via ;
        RECT 56.220 17.380 56.480 17.640 ;
        RECT 61.740 17.380 62.000 17.640 ;
      LAYER met2 ;
        RECT 61.800 17.670 61.940 54.000 ;
        RECT 56.220 17.350 56.480 17.670 ;
        RECT 61.740 17.350 62.000 17.670 ;
        RECT 56.280 2.400 56.420 17.350 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 80.110 16.900 80.430 16.960 ;
        RECT 82.410 16.900 82.730 16.960 ;
        RECT 80.110 16.760 82.730 16.900 ;
        RECT 80.110 16.700 80.430 16.760 ;
        RECT 82.410 16.700 82.730 16.760 ;
      LAYER via ;
        RECT 80.140 16.700 80.400 16.960 ;
        RECT 82.440 16.700 82.700 16.960 ;
      LAYER met2 ;
        RECT 82.500 16.990 82.640 54.000 ;
        RECT 80.140 16.670 80.400 16.990 ;
        RECT 82.440 16.670 82.700 16.990 ;
        RECT 80.200 2.400 80.340 16.670 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 103.570 17.920 103.890 17.980 ;
        RECT 109.550 17.920 109.870 17.980 ;
        RECT 103.570 17.780 109.870 17.920 ;
        RECT 103.570 17.720 103.890 17.780 ;
        RECT 109.550 17.720 109.870 17.780 ;
      LAYER via ;
        RECT 103.600 17.720 103.860 17.980 ;
        RECT 109.580 17.720 109.840 17.980 ;
      LAYER met2 ;
        RECT 109.640 18.010 109.780 54.000 ;
        RECT 103.600 17.690 103.860 18.010 ;
        RECT 109.580 17.690 109.840 18.010 ;
        RECT 103.660 2.400 103.800 17.690 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 127.490 17.580 127.810 17.640 ;
        RECT 130.710 17.580 131.030 17.640 ;
        RECT 127.490 17.440 131.030 17.580 ;
        RECT 127.490 17.380 127.810 17.440 ;
        RECT 130.710 17.380 131.030 17.440 ;
      LAYER via ;
        RECT 127.520 17.380 127.780 17.640 ;
        RECT 130.740 17.380 131.000 17.640 ;
      LAYER met2 ;
        RECT 130.800 17.670 130.940 54.000 ;
        RECT 127.520 17.350 127.780 17.670 ;
        RECT 130.740 17.350 131.000 17.670 ;
        RECT 127.580 2.400 127.720 17.350 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 27.210 372.880 27.530 372.940 ;
        RECT 27.210 372.740 54.000 372.880 ;
        RECT 27.210 372.680 27.530 372.740 ;
        RECT 26.290 2.960 26.610 3.020 ;
        RECT 27.210 2.960 27.530 3.020 ;
        RECT 26.290 2.820 27.530 2.960 ;
        RECT 26.290 2.760 26.610 2.820 ;
        RECT 27.210 2.760 27.530 2.820 ;
      LAYER via ;
        RECT 27.240 372.680 27.500 372.940 ;
        RECT 26.320 2.760 26.580 3.020 ;
        RECT 27.240 2.760 27.500 3.020 ;
      LAYER met2 ;
        RECT 27.240 372.650 27.500 372.970 ;
        RECT 27.300 3.050 27.440 372.650 ;
        RECT 26.320 2.730 26.580 3.050 ;
        RECT 27.240 2.730 27.500 3.050 ;
        RECT 26.380 2.400 26.520 2.730 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 34.110 386.480 34.430 386.540 ;
        RECT 34.110 386.340 54.000 386.480 ;
        RECT 34.110 386.280 34.430 386.340 ;
      LAYER via ;
        RECT 34.140 386.280 34.400 386.540 ;
      LAYER met2 ;
        RECT 34.140 386.250 34.400 386.570 ;
        RECT 34.200 3.130 34.340 386.250 ;
        RECT 32.360 2.990 34.340 3.130 ;
        RECT 32.360 2.400 32.500 2.990 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 653.730 14.180 654.050 14.240 ;
        RECT 656.950 14.180 657.270 14.240 ;
        RECT 674.430 14.180 674.750 14.240 ;
        RECT 692.370 14.180 692.690 14.240 ;
        RECT 710.310 14.180 710.630 14.240 ;
        RECT 728.250 14.180 728.570 14.240 ;
        RECT 746.190 14.180 746.510 14.240 ;
        RECT 763.670 14.180 763.990 14.240 ;
        RECT 781.610 14.180 781.930 14.240 ;
        RECT 799.550 14.180 799.870 14.240 ;
        RECT 817.490 14.180 817.810 14.240 ;
        RECT 835.430 14.180 835.750 14.240 ;
        RECT 852.910 14.180 853.230 14.240 ;
        RECT 870.850 14.180 871.170 14.240 ;
        RECT 888.790 14.180 889.110 14.240 ;
        RECT 906.730 14.180 907.050 14.240 ;
        RECT 924.210 14.180 924.530 14.240 ;
        RECT 942.150 14.180 942.470 14.240 ;
        RECT 960.090 14.180 960.410 14.240 ;
        RECT 978.030 14.180 978.350 14.240 ;
        RECT 995.970 14.180 996.290 14.240 ;
        RECT 1013.450 14.180 1013.770 14.240 ;
        RECT 1031.390 14.180 1031.710 14.240 ;
        RECT 1049.330 14.180 1049.650 14.240 ;
        RECT 1067.270 14.180 1067.590 14.240 ;
        RECT 1085.210 14.180 1085.530 14.240 ;
        RECT 1102.690 14.180 1103.010 14.240 ;
        RECT 1120.630 14.180 1120.950 14.240 ;
        RECT 1138.570 14.180 1138.890 14.240 ;
        RECT 1156.510 14.180 1156.830 14.240 ;
        RECT 1173.990 14.180 1174.310 14.240 ;
        RECT 1191.930 14.180 1192.250 14.240 ;
        RECT 1209.870 14.180 1210.190 14.240 ;
        RECT 1227.810 14.180 1228.130 14.240 ;
        RECT 1245.750 14.180 1246.070 14.240 ;
        RECT 1263.230 14.180 1263.550 14.240 ;
        RECT 1281.170 14.180 1281.490 14.240 ;
        RECT 1299.110 14.180 1299.430 14.240 ;
        RECT 1317.050 14.180 1317.370 14.240 ;
        RECT 1334.990 14.180 1335.310 14.240 ;
        RECT 1352.470 14.180 1352.790 14.240 ;
        RECT 1370.410 14.180 1370.730 14.240 ;
        RECT 1388.350 14.180 1388.670 14.240 ;
        RECT 1406.290 14.180 1406.610 14.240 ;
        RECT 1423.770 14.180 1424.090 14.240 ;
        RECT 1441.710 14.180 1442.030 14.240 ;
        RECT 1459.650 14.180 1459.970 14.240 ;
        RECT 1477.590 14.180 1477.910 14.240 ;
        RECT 1495.530 14.180 1495.850 14.240 ;
        RECT 1513.010 14.180 1513.330 14.240 ;
        RECT 1530.950 14.180 1531.270 14.240 ;
        RECT 1548.890 14.180 1549.210 14.240 ;
        RECT 1566.830 14.180 1567.150 14.240 ;
        RECT 1584.770 14.180 1585.090 14.240 ;
        RECT 1602.250 14.180 1602.570 14.240 ;
        RECT 1620.190 14.180 1620.510 14.240 ;
        RECT 1638.130 14.180 1638.450 14.240 ;
        RECT 1656.070 14.180 1656.390 14.240 ;
        RECT 1673.550 14.180 1673.870 14.240 ;
        RECT 1691.490 14.180 1691.810 14.240 ;
        RECT 1709.430 14.180 1709.750 14.240 ;
        RECT 1727.370 14.180 1727.690 14.240 ;
        RECT 1745.310 14.180 1745.630 14.240 ;
        RECT 1762.790 14.180 1763.110 14.240 ;
        RECT 1780.730 14.180 1781.050 14.240 ;
        RECT 1798.670 14.180 1798.990 14.240 ;
        RECT 1816.610 14.180 1816.930 14.240 ;
        RECT 1834.550 14.180 1834.870 14.240 ;
        RECT 1852.030 14.180 1852.350 14.240 ;
        RECT 1869.970 14.180 1870.290 14.240 ;
        RECT 1887.910 14.180 1888.230 14.240 ;
        RECT 1905.850 14.180 1906.170 14.240 ;
        RECT 1923.330 14.180 1923.650 14.240 ;
        RECT 1941.270 14.180 1941.590 14.240 ;
        RECT 1959.210 14.180 1959.530 14.240 ;
        RECT 1977.150 14.180 1977.470 14.240 ;
        RECT 1995.090 14.180 1995.410 14.240 ;
        RECT 2012.570 14.180 2012.890 14.240 ;
        RECT 2030.510 14.180 2030.830 14.240 ;
        RECT 2048.450 14.180 2048.770 14.240 ;
        RECT 2066.390 14.180 2066.710 14.240 ;
        RECT 2084.330 14.180 2084.650 14.240 ;
        RECT 2101.810 14.180 2102.130 14.240 ;
        RECT 2119.750 14.180 2120.070 14.240 ;
        RECT 2137.690 14.180 2138.010 14.240 ;
        RECT 2155.630 14.180 2155.950 14.240 ;
        RECT 2173.110 14.180 2173.430 14.240 ;
        RECT 2191.050 14.180 2191.370 14.240 ;
        RECT 2208.990 14.180 2209.310 14.240 ;
        RECT 2226.930 14.180 2227.250 14.240 ;
        RECT 2244.870 14.180 2245.190 14.240 ;
        RECT 2262.350 14.180 2262.670 14.240 ;
        RECT 2280.290 14.180 2280.610 14.240 ;
        RECT 2298.230 14.180 2298.550 14.240 ;
        RECT 2316.170 14.180 2316.490 14.240 ;
        RECT 2334.110 14.180 2334.430 14.240 ;
        RECT 2351.590 14.180 2351.910 14.240 ;
        RECT 2369.530 14.180 2369.850 14.240 ;
        RECT 2387.470 14.180 2387.790 14.240 ;
        RECT 2405.410 14.180 2405.730 14.240 ;
        RECT 2422.890 14.180 2423.210 14.240 ;
        RECT 2440.830 14.180 2441.150 14.240 ;
        RECT 2458.770 14.180 2459.090 14.240 ;
        RECT 2476.710 14.180 2477.030 14.240 ;
        RECT 2494.650 14.180 2494.970 14.240 ;
        RECT 2512.130 14.180 2512.450 14.240 ;
        RECT 2530.070 14.180 2530.390 14.240 ;
        RECT 2548.010 14.180 2548.330 14.240 ;
        RECT 2565.950 14.180 2566.270 14.240 ;
        RECT 2583.890 14.180 2584.210 14.240 ;
        RECT 2601.370 14.180 2601.690 14.240 ;
        RECT 2619.310 14.180 2619.630 14.240 ;
        RECT 2637.250 14.180 2637.570 14.240 ;
        RECT 2655.190 14.180 2655.510 14.240 ;
        RECT 2672.670 14.180 2672.990 14.240 ;
        RECT 2690.610 14.180 2690.930 14.240 ;
        RECT 2708.550 14.180 2708.870 14.240 ;
        RECT 2726.490 14.180 2726.810 14.240 ;
        RECT 2744.430 14.180 2744.750 14.240 ;
        RECT 2761.910 14.180 2762.230 14.240 ;
        RECT 2779.850 14.180 2780.170 14.240 ;
        RECT 2797.790 14.180 2798.110 14.240 ;
        RECT 2815.730 14.180 2816.050 14.240 ;
        RECT 2833.670 14.180 2833.990 14.240 ;
        RECT 2851.150 14.180 2851.470 14.240 ;
        RECT 2869.090 14.180 2869.410 14.240 ;
        RECT 2887.030 14.180 2887.350 14.240 ;
        RECT 2904.970 14.180 2905.290 14.240 ;
        RECT 653.730 14.040 2905.290 14.180 ;
        RECT 653.730 13.980 654.050 14.040 ;
        RECT 656.950 13.980 657.270 14.040 ;
        RECT 674.430 13.980 674.750 14.040 ;
        RECT 692.370 13.980 692.690 14.040 ;
        RECT 710.310 13.980 710.630 14.040 ;
        RECT 728.250 13.980 728.570 14.040 ;
        RECT 746.190 13.980 746.510 14.040 ;
        RECT 763.670 13.980 763.990 14.040 ;
        RECT 781.610 13.980 781.930 14.040 ;
        RECT 799.550 13.980 799.870 14.040 ;
        RECT 817.490 13.980 817.810 14.040 ;
        RECT 835.430 13.980 835.750 14.040 ;
        RECT 852.910 13.980 853.230 14.040 ;
        RECT 870.850 13.980 871.170 14.040 ;
        RECT 888.790 13.980 889.110 14.040 ;
        RECT 906.730 13.980 907.050 14.040 ;
        RECT 924.210 13.980 924.530 14.040 ;
        RECT 942.150 13.980 942.470 14.040 ;
        RECT 960.090 13.980 960.410 14.040 ;
        RECT 978.030 13.980 978.350 14.040 ;
        RECT 995.970 13.980 996.290 14.040 ;
        RECT 1013.450 13.980 1013.770 14.040 ;
        RECT 1031.390 13.980 1031.710 14.040 ;
        RECT 1049.330 13.980 1049.650 14.040 ;
        RECT 1067.270 13.980 1067.590 14.040 ;
        RECT 1085.210 13.980 1085.530 14.040 ;
        RECT 1102.690 13.980 1103.010 14.040 ;
        RECT 1120.630 13.980 1120.950 14.040 ;
        RECT 1138.570 13.980 1138.890 14.040 ;
        RECT 1156.510 13.980 1156.830 14.040 ;
        RECT 1173.990 13.980 1174.310 14.040 ;
        RECT 1191.930 13.980 1192.250 14.040 ;
        RECT 1209.870 13.980 1210.190 14.040 ;
        RECT 1227.810 13.980 1228.130 14.040 ;
        RECT 1245.750 13.980 1246.070 14.040 ;
        RECT 1263.230 13.980 1263.550 14.040 ;
        RECT 1281.170 13.980 1281.490 14.040 ;
        RECT 1299.110 13.980 1299.430 14.040 ;
        RECT 1317.050 13.980 1317.370 14.040 ;
        RECT 1334.990 13.980 1335.310 14.040 ;
        RECT 1352.470 13.980 1352.790 14.040 ;
        RECT 1370.410 13.980 1370.730 14.040 ;
        RECT 1388.350 13.980 1388.670 14.040 ;
        RECT 1406.290 13.980 1406.610 14.040 ;
        RECT 1423.770 13.980 1424.090 14.040 ;
        RECT 1441.710 13.980 1442.030 14.040 ;
        RECT 1459.650 13.980 1459.970 14.040 ;
        RECT 1477.590 13.980 1477.910 14.040 ;
        RECT 1495.530 13.980 1495.850 14.040 ;
        RECT 1513.010 13.980 1513.330 14.040 ;
        RECT 1530.950 13.980 1531.270 14.040 ;
        RECT 1548.890 13.980 1549.210 14.040 ;
        RECT 1566.830 13.980 1567.150 14.040 ;
        RECT 1584.770 13.980 1585.090 14.040 ;
        RECT 1602.250 13.980 1602.570 14.040 ;
        RECT 1620.190 13.980 1620.510 14.040 ;
        RECT 1638.130 13.980 1638.450 14.040 ;
        RECT 1656.070 13.980 1656.390 14.040 ;
        RECT 1673.550 13.980 1673.870 14.040 ;
        RECT 1691.490 13.980 1691.810 14.040 ;
        RECT 1709.430 13.980 1709.750 14.040 ;
        RECT 1727.370 13.980 1727.690 14.040 ;
        RECT 1745.310 13.980 1745.630 14.040 ;
        RECT 1762.790 13.980 1763.110 14.040 ;
        RECT 1780.730 13.980 1781.050 14.040 ;
        RECT 1798.670 13.980 1798.990 14.040 ;
        RECT 1816.610 13.980 1816.930 14.040 ;
        RECT 1834.550 13.980 1834.870 14.040 ;
        RECT 1852.030 13.980 1852.350 14.040 ;
        RECT 1869.970 13.980 1870.290 14.040 ;
        RECT 1887.910 13.980 1888.230 14.040 ;
        RECT 1905.850 13.980 1906.170 14.040 ;
        RECT 1923.330 13.980 1923.650 14.040 ;
        RECT 1941.270 13.980 1941.590 14.040 ;
        RECT 1959.210 13.980 1959.530 14.040 ;
        RECT 1977.150 13.980 1977.470 14.040 ;
        RECT 1995.090 13.980 1995.410 14.040 ;
        RECT 2012.570 13.980 2012.890 14.040 ;
        RECT 2030.510 13.980 2030.830 14.040 ;
        RECT 2048.450 13.980 2048.770 14.040 ;
        RECT 2066.390 13.980 2066.710 14.040 ;
        RECT 2084.330 13.980 2084.650 14.040 ;
        RECT 2101.810 13.980 2102.130 14.040 ;
        RECT 2119.750 13.980 2120.070 14.040 ;
        RECT 2137.690 13.980 2138.010 14.040 ;
        RECT 2155.630 13.980 2155.950 14.040 ;
        RECT 2173.110 13.980 2173.430 14.040 ;
        RECT 2191.050 13.980 2191.370 14.040 ;
        RECT 2208.990 13.980 2209.310 14.040 ;
        RECT 2226.930 13.980 2227.250 14.040 ;
        RECT 2244.870 13.980 2245.190 14.040 ;
        RECT 2262.350 13.980 2262.670 14.040 ;
        RECT 2280.290 13.980 2280.610 14.040 ;
        RECT 2298.230 13.980 2298.550 14.040 ;
        RECT 2316.170 13.980 2316.490 14.040 ;
        RECT 2334.110 13.980 2334.430 14.040 ;
        RECT 2351.590 13.980 2351.910 14.040 ;
        RECT 2369.530 13.980 2369.850 14.040 ;
        RECT 2387.470 13.980 2387.790 14.040 ;
        RECT 2405.410 13.980 2405.730 14.040 ;
        RECT 2422.890 13.980 2423.210 14.040 ;
        RECT 2440.830 13.980 2441.150 14.040 ;
        RECT 2458.770 13.980 2459.090 14.040 ;
        RECT 2476.710 13.980 2477.030 14.040 ;
        RECT 2494.650 13.980 2494.970 14.040 ;
        RECT 2512.130 13.980 2512.450 14.040 ;
        RECT 2530.070 13.980 2530.390 14.040 ;
        RECT 2548.010 13.980 2548.330 14.040 ;
        RECT 2565.950 13.980 2566.270 14.040 ;
        RECT 2583.890 13.980 2584.210 14.040 ;
        RECT 2601.370 13.980 2601.690 14.040 ;
        RECT 2619.310 13.980 2619.630 14.040 ;
        RECT 2637.250 13.980 2637.570 14.040 ;
        RECT 2655.190 13.980 2655.510 14.040 ;
        RECT 2672.670 13.980 2672.990 14.040 ;
        RECT 2690.610 13.980 2690.930 14.040 ;
        RECT 2708.550 13.980 2708.870 14.040 ;
        RECT 2726.490 13.980 2726.810 14.040 ;
        RECT 2744.430 13.980 2744.750 14.040 ;
        RECT 2761.910 13.980 2762.230 14.040 ;
        RECT 2779.850 13.980 2780.170 14.040 ;
        RECT 2797.790 13.980 2798.110 14.040 ;
        RECT 2815.730 13.980 2816.050 14.040 ;
        RECT 2833.670 13.980 2833.990 14.040 ;
        RECT 2851.150 13.980 2851.470 14.040 ;
        RECT 2869.090 13.980 2869.410 14.040 ;
        RECT 2887.030 13.980 2887.350 14.040 ;
        RECT 2904.970 13.980 2905.290 14.040 ;
        RECT 639.010 2.960 639.330 3.020 ;
        RECT 656.950 2.960 657.270 3.020 ;
        RECT 639.010 2.820 657.270 2.960 ;
        RECT 639.010 2.760 639.330 2.820 ;
        RECT 656.950 2.760 657.270 2.820 ;
      LAYER via ;
        RECT 653.760 13.980 654.020 14.240 ;
        RECT 656.980 13.980 657.240 14.240 ;
        RECT 674.460 13.980 674.720 14.240 ;
        RECT 692.400 13.980 692.660 14.240 ;
        RECT 710.340 13.980 710.600 14.240 ;
        RECT 728.280 13.980 728.540 14.240 ;
        RECT 746.220 13.980 746.480 14.240 ;
        RECT 763.700 13.980 763.960 14.240 ;
        RECT 781.640 13.980 781.900 14.240 ;
        RECT 799.580 13.980 799.840 14.240 ;
        RECT 817.520 13.980 817.780 14.240 ;
        RECT 835.460 13.980 835.720 14.240 ;
        RECT 852.940 13.980 853.200 14.240 ;
        RECT 870.880 13.980 871.140 14.240 ;
        RECT 888.820 13.980 889.080 14.240 ;
        RECT 906.760 13.980 907.020 14.240 ;
        RECT 924.240 13.980 924.500 14.240 ;
        RECT 942.180 13.980 942.440 14.240 ;
        RECT 960.120 13.980 960.380 14.240 ;
        RECT 978.060 13.980 978.320 14.240 ;
        RECT 996.000 13.980 996.260 14.240 ;
        RECT 1013.480 13.980 1013.740 14.240 ;
        RECT 1031.420 13.980 1031.680 14.240 ;
        RECT 1049.360 13.980 1049.620 14.240 ;
        RECT 1067.300 13.980 1067.560 14.240 ;
        RECT 1085.240 13.980 1085.500 14.240 ;
        RECT 1102.720 13.980 1102.980 14.240 ;
        RECT 1120.660 13.980 1120.920 14.240 ;
        RECT 1138.600 13.980 1138.860 14.240 ;
        RECT 1156.540 13.980 1156.800 14.240 ;
        RECT 1174.020 13.980 1174.280 14.240 ;
        RECT 1191.960 13.980 1192.220 14.240 ;
        RECT 1209.900 13.980 1210.160 14.240 ;
        RECT 1227.840 13.980 1228.100 14.240 ;
        RECT 1245.780 13.980 1246.040 14.240 ;
        RECT 1263.260 13.980 1263.520 14.240 ;
        RECT 1281.200 13.980 1281.460 14.240 ;
        RECT 1299.140 13.980 1299.400 14.240 ;
        RECT 1317.080 13.980 1317.340 14.240 ;
        RECT 1335.020 13.980 1335.280 14.240 ;
        RECT 1352.500 13.980 1352.760 14.240 ;
        RECT 1370.440 13.980 1370.700 14.240 ;
        RECT 1388.380 13.980 1388.640 14.240 ;
        RECT 1406.320 13.980 1406.580 14.240 ;
        RECT 1423.800 13.980 1424.060 14.240 ;
        RECT 1441.740 13.980 1442.000 14.240 ;
        RECT 1459.680 13.980 1459.940 14.240 ;
        RECT 1477.620 13.980 1477.880 14.240 ;
        RECT 1495.560 13.980 1495.820 14.240 ;
        RECT 1513.040 13.980 1513.300 14.240 ;
        RECT 1530.980 13.980 1531.240 14.240 ;
        RECT 1548.920 13.980 1549.180 14.240 ;
        RECT 1566.860 13.980 1567.120 14.240 ;
        RECT 1584.800 13.980 1585.060 14.240 ;
        RECT 1602.280 13.980 1602.540 14.240 ;
        RECT 1620.220 13.980 1620.480 14.240 ;
        RECT 1638.160 13.980 1638.420 14.240 ;
        RECT 1656.100 13.980 1656.360 14.240 ;
        RECT 1673.580 13.980 1673.840 14.240 ;
        RECT 1691.520 13.980 1691.780 14.240 ;
        RECT 1709.460 13.980 1709.720 14.240 ;
        RECT 1727.400 13.980 1727.660 14.240 ;
        RECT 1745.340 13.980 1745.600 14.240 ;
        RECT 1762.820 13.980 1763.080 14.240 ;
        RECT 1780.760 13.980 1781.020 14.240 ;
        RECT 1798.700 13.980 1798.960 14.240 ;
        RECT 1816.640 13.980 1816.900 14.240 ;
        RECT 1834.580 13.980 1834.840 14.240 ;
        RECT 1852.060 13.980 1852.320 14.240 ;
        RECT 1870.000 13.980 1870.260 14.240 ;
        RECT 1887.940 13.980 1888.200 14.240 ;
        RECT 1905.880 13.980 1906.140 14.240 ;
        RECT 1923.360 13.980 1923.620 14.240 ;
        RECT 1941.300 13.980 1941.560 14.240 ;
        RECT 1959.240 13.980 1959.500 14.240 ;
        RECT 1977.180 13.980 1977.440 14.240 ;
        RECT 1995.120 13.980 1995.380 14.240 ;
        RECT 2012.600 13.980 2012.860 14.240 ;
        RECT 2030.540 13.980 2030.800 14.240 ;
        RECT 2048.480 13.980 2048.740 14.240 ;
        RECT 2066.420 13.980 2066.680 14.240 ;
        RECT 2084.360 13.980 2084.620 14.240 ;
        RECT 2101.840 13.980 2102.100 14.240 ;
        RECT 2119.780 13.980 2120.040 14.240 ;
        RECT 2137.720 13.980 2137.980 14.240 ;
        RECT 2155.660 13.980 2155.920 14.240 ;
        RECT 2173.140 13.980 2173.400 14.240 ;
        RECT 2191.080 13.980 2191.340 14.240 ;
        RECT 2209.020 13.980 2209.280 14.240 ;
        RECT 2226.960 13.980 2227.220 14.240 ;
        RECT 2244.900 13.980 2245.160 14.240 ;
        RECT 2262.380 13.980 2262.640 14.240 ;
        RECT 2280.320 13.980 2280.580 14.240 ;
        RECT 2298.260 13.980 2298.520 14.240 ;
        RECT 2316.200 13.980 2316.460 14.240 ;
        RECT 2334.140 13.980 2334.400 14.240 ;
        RECT 2351.620 13.980 2351.880 14.240 ;
        RECT 2369.560 13.980 2369.820 14.240 ;
        RECT 2387.500 13.980 2387.760 14.240 ;
        RECT 2405.440 13.980 2405.700 14.240 ;
        RECT 2422.920 13.980 2423.180 14.240 ;
        RECT 2440.860 13.980 2441.120 14.240 ;
        RECT 2458.800 13.980 2459.060 14.240 ;
        RECT 2476.740 13.980 2477.000 14.240 ;
        RECT 2494.680 13.980 2494.940 14.240 ;
        RECT 2512.160 13.980 2512.420 14.240 ;
        RECT 2530.100 13.980 2530.360 14.240 ;
        RECT 2548.040 13.980 2548.300 14.240 ;
        RECT 2565.980 13.980 2566.240 14.240 ;
        RECT 2583.920 13.980 2584.180 14.240 ;
        RECT 2601.400 13.980 2601.660 14.240 ;
        RECT 2619.340 13.980 2619.600 14.240 ;
        RECT 2637.280 13.980 2637.540 14.240 ;
        RECT 2655.220 13.980 2655.480 14.240 ;
        RECT 2672.700 13.980 2672.960 14.240 ;
        RECT 2690.640 13.980 2690.900 14.240 ;
        RECT 2708.580 13.980 2708.840 14.240 ;
        RECT 2726.520 13.980 2726.780 14.240 ;
        RECT 2744.460 13.980 2744.720 14.240 ;
        RECT 2761.940 13.980 2762.200 14.240 ;
        RECT 2779.880 13.980 2780.140 14.240 ;
        RECT 2797.820 13.980 2798.080 14.240 ;
        RECT 2815.760 13.980 2816.020 14.240 ;
        RECT 2833.700 13.980 2833.960 14.240 ;
        RECT 2851.180 13.980 2851.440 14.240 ;
        RECT 2869.120 13.980 2869.380 14.240 ;
        RECT 2887.060 13.980 2887.320 14.240 ;
        RECT 2905.000 13.980 2905.260 14.240 ;
        RECT 639.040 2.760 639.300 3.020 ;
        RECT 656.980 2.760 657.240 3.020 ;
      LAYER met2 ;
        RECT 653.820 14.270 653.960 54.000 ;
        RECT 653.760 13.950 654.020 14.270 ;
        RECT 656.980 13.950 657.240 14.270 ;
        RECT 674.460 13.950 674.720 14.270 ;
        RECT 692.400 13.950 692.660 14.270 ;
        RECT 710.340 13.950 710.600 14.270 ;
        RECT 728.280 13.950 728.540 14.270 ;
        RECT 746.220 13.950 746.480 14.270 ;
        RECT 763.700 13.950 763.960 14.270 ;
        RECT 781.640 13.950 781.900 14.270 ;
        RECT 799.580 13.950 799.840 14.270 ;
        RECT 817.520 13.950 817.780 14.270 ;
        RECT 835.460 13.950 835.720 14.270 ;
        RECT 852.940 13.950 853.200 14.270 ;
        RECT 870.880 13.950 871.140 14.270 ;
        RECT 888.820 13.950 889.080 14.270 ;
        RECT 906.760 13.950 907.020 14.270 ;
        RECT 924.240 13.950 924.500 14.270 ;
        RECT 942.180 13.950 942.440 14.270 ;
        RECT 960.120 13.950 960.380 14.270 ;
        RECT 978.060 13.950 978.320 14.270 ;
        RECT 996.000 13.950 996.260 14.270 ;
        RECT 1013.480 13.950 1013.740 14.270 ;
        RECT 1031.420 13.950 1031.680 14.270 ;
        RECT 1049.360 13.950 1049.620 14.270 ;
        RECT 1067.300 13.950 1067.560 14.270 ;
        RECT 1085.240 13.950 1085.500 14.270 ;
        RECT 1102.720 13.950 1102.980 14.270 ;
        RECT 1120.660 13.950 1120.920 14.270 ;
        RECT 1138.600 13.950 1138.860 14.270 ;
        RECT 1156.540 13.950 1156.800 14.270 ;
        RECT 1174.020 13.950 1174.280 14.270 ;
        RECT 1191.960 13.950 1192.220 14.270 ;
        RECT 1209.900 13.950 1210.160 14.270 ;
        RECT 1227.840 13.950 1228.100 14.270 ;
        RECT 1245.780 13.950 1246.040 14.270 ;
        RECT 1263.260 13.950 1263.520 14.270 ;
        RECT 1281.200 13.950 1281.460 14.270 ;
        RECT 1299.140 13.950 1299.400 14.270 ;
        RECT 1317.080 13.950 1317.340 14.270 ;
        RECT 1335.020 13.950 1335.280 14.270 ;
        RECT 1352.500 13.950 1352.760 14.270 ;
        RECT 1370.440 13.950 1370.700 14.270 ;
        RECT 1388.380 13.950 1388.640 14.270 ;
        RECT 1406.320 13.950 1406.580 14.270 ;
        RECT 1423.800 13.950 1424.060 14.270 ;
        RECT 1441.740 13.950 1442.000 14.270 ;
        RECT 1459.680 13.950 1459.940 14.270 ;
        RECT 1477.620 13.950 1477.880 14.270 ;
        RECT 1495.560 13.950 1495.820 14.270 ;
        RECT 1513.040 13.950 1513.300 14.270 ;
        RECT 1530.980 13.950 1531.240 14.270 ;
        RECT 1548.920 13.950 1549.180 14.270 ;
        RECT 1566.860 13.950 1567.120 14.270 ;
        RECT 1584.800 13.950 1585.060 14.270 ;
        RECT 1602.280 13.950 1602.540 14.270 ;
        RECT 1620.220 13.950 1620.480 14.270 ;
        RECT 1638.160 13.950 1638.420 14.270 ;
        RECT 1656.100 13.950 1656.360 14.270 ;
        RECT 1673.580 13.950 1673.840 14.270 ;
        RECT 1691.520 13.950 1691.780 14.270 ;
        RECT 1709.460 13.950 1709.720 14.270 ;
        RECT 1727.400 13.950 1727.660 14.270 ;
        RECT 1745.340 13.950 1745.600 14.270 ;
        RECT 1762.820 13.950 1763.080 14.270 ;
        RECT 1780.760 13.950 1781.020 14.270 ;
        RECT 1798.700 13.950 1798.960 14.270 ;
        RECT 1816.640 13.950 1816.900 14.270 ;
        RECT 1834.580 13.950 1834.840 14.270 ;
        RECT 1852.060 13.950 1852.320 14.270 ;
        RECT 1870.000 13.950 1870.260 14.270 ;
        RECT 1887.940 13.950 1888.200 14.270 ;
        RECT 1905.880 13.950 1906.140 14.270 ;
        RECT 1923.360 13.950 1923.620 14.270 ;
        RECT 1941.300 13.950 1941.560 14.270 ;
        RECT 1959.240 13.950 1959.500 14.270 ;
        RECT 1977.180 13.950 1977.440 14.270 ;
        RECT 1995.120 13.950 1995.380 14.270 ;
        RECT 2012.600 13.950 2012.860 14.270 ;
        RECT 2030.540 13.950 2030.800 14.270 ;
        RECT 2048.480 13.950 2048.740 14.270 ;
        RECT 2066.420 13.950 2066.680 14.270 ;
        RECT 2084.360 13.950 2084.620 14.270 ;
        RECT 2101.840 13.950 2102.100 14.270 ;
        RECT 2119.780 13.950 2120.040 14.270 ;
        RECT 2137.720 13.950 2137.980 14.270 ;
        RECT 2155.660 13.950 2155.920 14.270 ;
        RECT 2173.140 13.950 2173.400 14.270 ;
        RECT 2191.080 13.950 2191.340 14.270 ;
        RECT 2209.020 13.950 2209.280 14.270 ;
        RECT 2226.960 13.950 2227.220 14.270 ;
        RECT 2244.900 13.950 2245.160 14.270 ;
        RECT 2262.380 13.950 2262.640 14.270 ;
        RECT 2280.320 13.950 2280.580 14.270 ;
        RECT 2298.260 13.950 2298.520 14.270 ;
        RECT 2316.200 13.950 2316.460 14.270 ;
        RECT 2334.140 13.950 2334.400 14.270 ;
        RECT 2351.620 13.950 2351.880 14.270 ;
        RECT 2369.560 13.950 2369.820 14.270 ;
        RECT 2387.500 13.950 2387.760 14.270 ;
        RECT 2405.440 13.950 2405.700 14.270 ;
        RECT 2422.920 13.950 2423.180 14.270 ;
        RECT 2440.860 13.950 2441.120 14.270 ;
        RECT 2458.800 13.950 2459.060 14.270 ;
        RECT 2476.740 13.950 2477.000 14.270 ;
        RECT 2494.680 13.950 2494.940 14.270 ;
        RECT 2512.160 13.950 2512.420 14.270 ;
        RECT 2530.100 13.950 2530.360 14.270 ;
        RECT 2548.040 13.950 2548.300 14.270 ;
        RECT 2565.980 13.950 2566.240 14.270 ;
        RECT 2583.920 13.950 2584.180 14.270 ;
        RECT 2601.400 13.950 2601.660 14.270 ;
        RECT 2619.340 13.950 2619.600 14.270 ;
        RECT 2637.280 13.950 2637.540 14.270 ;
        RECT 2655.220 13.950 2655.480 14.270 ;
        RECT 2672.700 13.950 2672.960 14.270 ;
        RECT 2690.640 13.950 2690.900 14.270 ;
        RECT 2708.580 13.950 2708.840 14.270 ;
        RECT 2726.520 13.950 2726.780 14.270 ;
        RECT 2744.460 13.950 2744.720 14.270 ;
        RECT 2761.940 13.950 2762.200 14.270 ;
        RECT 2779.880 13.950 2780.140 14.270 ;
        RECT 2797.820 13.950 2798.080 14.270 ;
        RECT 2815.760 13.950 2816.020 14.270 ;
        RECT 2833.700 13.950 2833.960 14.270 ;
        RECT 2851.180 13.950 2851.440 14.270 ;
        RECT 2869.120 13.950 2869.380 14.270 ;
        RECT 2887.060 13.950 2887.320 14.270 ;
        RECT 2905.000 13.950 2905.260 14.270 ;
        RECT 657.040 3.050 657.180 13.950 ;
        RECT 639.040 2.730 639.300 3.050 ;
        RECT 656.980 2.730 657.240 3.050 ;
        RECT 639.100 2.400 639.240 2.730 ;
        RECT 657.040 2.400 657.180 2.730 ;
        RECT 674.520 2.400 674.660 13.950 ;
        RECT 692.460 2.400 692.600 13.950 ;
        RECT 710.400 2.400 710.540 13.950 ;
        RECT 728.340 2.400 728.480 13.950 ;
        RECT 746.280 2.400 746.420 13.950 ;
        RECT 763.760 2.400 763.900 13.950 ;
        RECT 781.700 2.400 781.840 13.950 ;
        RECT 799.640 2.400 799.780 13.950 ;
        RECT 817.580 2.400 817.720 13.950 ;
        RECT 835.520 2.400 835.660 13.950 ;
        RECT 853.000 2.400 853.140 13.950 ;
        RECT 870.940 2.400 871.080 13.950 ;
        RECT 888.880 2.400 889.020 13.950 ;
        RECT 906.820 2.400 906.960 13.950 ;
        RECT 924.300 2.400 924.440 13.950 ;
        RECT 942.240 2.400 942.380 13.950 ;
        RECT 960.180 2.400 960.320 13.950 ;
        RECT 978.120 2.400 978.260 13.950 ;
        RECT 996.060 2.400 996.200 13.950 ;
        RECT 1013.540 2.400 1013.680 13.950 ;
        RECT 1031.480 2.400 1031.620 13.950 ;
        RECT 1049.420 2.400 1049.560 13.950 ;
        RECT 1067.360 2.400 1067.500 13.950 ;
        RECT 1085.300 2.400 1085.440 13.950 ;
        RECT 1102.780 2.400 1102.920 13.950 ;
        RECT 1120.720 2.400 1120.860 13.950 ;
        RECT 1138.660 2.400 1138.800 13.950 ;
        RECT 1156.600 2.400 1156.740 13.950 ;
        RECT 1174.080 2.400 1174.220 13.950 ;
        RECT 1192.020 2.400 1192.160 13.950 ;
        RECT 1209.960 2.400 1210.100 13.950 ;
        RECT 1227.900 2.400 1228.040 13.950 ;
        RECT 1245.840 2.400 1245.980 13.950 ;
        RECT 1263.320 2.400 1263.460 13.950 ;
        RECT 1281.260 2.400 1281.400 13.950 ;
        RECT 1299.200 2.400 1299.340 13.950 ;
        RECT 1317.140 2.400 1317.280 13.950 ;
        RECT 1335.080 2.400 1335.220 13.950 ;
        RECT 1352.560 2.400 1352.700 13.950 ;
        RECT 1370.500 2.400 1370.640 13.950 ;
        RECT 1388.440 2.400 1388.580 13.950 ;
        RECT 1406.380 2.400 1406.520 13.950 ;
        RECT 1423.860 2.400 1424.000 13.950 ;
        RECT 1441.800 2.400 1441.940 13.950 ;
        RECT 1459.740 2.400 1459.880 13.950 ;
        RECT 1477.680 2.400 1477.820 13.950 ;
        RECT 1495.620 2.400 1495.760 13.950 ;
        RECT 1513.100 2.400 1513.240 13.950 ;
        RECT 1531.040 2.400 1531.180 13.950 ;
        RECT 1548.980 2.400 1549.120 13.950 ;
        RECT 1566.920 2.400 1567.060 13.950 ;
        RECT 1584.860 2.400 1585.000 13.950 ;
        RECT 1602.340 2.400 1602.480 13.950 ;
        RECT 1620.280 2.400 1620.420 13.950 ;
        RECT 1638.220 2.400 1638.360 13.950 ;
        RECT 1656.160 2.400 1656.300 13.950 ;
        RECT 1673.640 2.400 1673.780 13.950 ;
        RECT 1691.580 2.400 1691.720 13.950 ;
        RECT 1709.520 2.400 1709.660 13.950 ;
        RECT 1727.460 2.400 1727.600 13.950 ;
        RECT 1745.400 2.400 1745.540 13.950 ;
        RECT 1762.880 2.400 1763.020 13.950 ;
        RECT 1780.820 2.400 1780.960 13.950 ;
        RECT 1798.760 2.400 1798.900 13.950 ;
        RECT 1816.700 2.400 1816.840 13.950 ;
        RECT 1834.640 2.400 1834.780 13.950 ;
        RECT 1852.120 2.400 1852.260 13.950 ;
        RECT 1870.060 2.400 1870.200 13.950 ;
        RECT 1888.000 2.400 1888.140 13.950 ;
        RECT 1905.940 2.400 1906.080 13.950 ;
        RECT 1923.420 2.400 1923.560 13.950 ;
        RECT 1941.360 2.400 1941.500 13.950 ;
        RECT 1959.300 2.400 1959.440 13.950 ;
        RECT 1977.240 2.400 1977.380 13.950 ;
        RECT 1995.180 2.400 1995.320 13.950 ;
        RECT 2012.660 2.400 2012.800 13.950 ;
        RECT 2030.600 2.400 2030.740 13.950 ;
        RECT 2048.540 2.400 2048.680 13.950 ;
        RECT 2066.480 2.400 2066.620 13.950 ;
        RECT 2084.420 2.400 2084.560 13.950 ;
        RECT 2101.900 2.400 2102.040 13.950 ;
        RECT 2119.840 2.400 2119.980 13.950 ;
        RECT 2137.780 2.400 2137.920 13.950 ;
        RECT 2155.720 2.400 2155.860 13.950 ;
        RECT 2173.200 2.400 2173.340 13.950 ;
        RECT 2191.140 2.400 2191.280 13.950 ;
        RECT 2209.080 2.400 2209.220 13.950 ;
        RECT 2227.020 2.400 2227.160 13.950 ;
        RECT 2244.960 2.400 2245.100 13.950 ;
        RECT 2262.440 2.400 2262.580 13.950 ;
        RECT 2280.380 2.400 2280.520 13.950 ;
        RECT 2298.320 2.400 2298.460 13.950 ;
        RECT 2316.260 2.400 2316.400 13.950 ;
        RECT 2334.200 2.400 2334.340 13.950 ;
        RECT 2351.680 2.400 2351.820 13.950 ;
        RECT 2369.620 2.400 2369.760 13.950 ;
        RECT 2387.560 2.400 2387.700 13.950 ;
        RECT 2405.500 2.400 2405.640 13.950 ;
        RECT 2422.980 2.400 2423.120 13.950 ;
        RECT 2440.920 2.400 2441.060 13.950 ;
        RECT 2458.860 2.400 2459.000 13.950 ;
        RECT 2476.800 2.400 2476.940 13.950 ;
        RECT 2494.740 2.400 2494.880 13.950 ;
        RECT 2512.220 2.400 2512.360 13.950 ;
        RECT 2530.160 2.400 2530.300 13.950 ;
        RECT 2548.100 2.400 2548.240 13.950 ;
        RECT 2566.040 2.400 2566.180 13.950 ;
        RECT 2583.980 2.400 2584.120 13.950 ;
        RECT 2601.460 2.400 2601.600 13.950 ;
        RECT 2619.400 2.400 2619.540 13.950 ;
        RECT 2637.340 2.400 2637.480 13.950 ;
        RECT 2655.280 2.400 2655.420 13.950 ;
        RECT 2672.760 2.400 2672.900 13.950 ;
        RECT 2690.700 2.400 2690.840 13.950 ;
        RECT 2708.640 2.400 2708.780 13.950 ;
        RECT 2726.580 2.400 2726.720 13.950 ;
        RECT 2744.520 2.400 2744.660 13.950 ;
        RECT 2762.000 2.400 2762.140 13.950 ;
        RECT 2779.940 2.400 2780.080 13.950 ;
        RECT 2797.880 2.400 2798.020 13.950 ;
        RECT 2815.820 2.400 2815.960 13.950 ;
        RECT 2833.760 2.400 2833.900 13.950 ;
        RECT 2851.240 2.400 2851.380 13.950 ;
        RECT 2869.180 2.400 2869.320 13.950 ;
        RECT 2887.120 2.400 2887.260 13.950 ;
        RECT 2905.060 2.400 2905.200 13.950 ;
        RECT 638.890 -4.800 639.450 2.400 ;
        RECT 656.830 -4.800 657.390 2.400 ;
        RECT 674.310 -4.800 674.870 2.400 ;
        RECT 692.250 -4.800 692.810 2.400 ;
        RECT 710.190 -4.800 710.750 2.400 ;
        RECT 728.130 -4.800 728.690 2.400 ;
        RECT 746.070 -4.800 746.630 2.400 ;
        RECT 763.550 -4.800 764.110 2.400 ;
        RECT 781.490 -4.800 782.050 2.400 ;
        RECT 799.430 -4.800 799.990 2.400 ;
        RECT 817.370 -4.800 817.930 2.400 ;
        RECT 835.310 -4.800 835.870 2.400 ;
        RECT 852.790 -4.800 853.350 2.400 ;
        RECT 870.730 -4.800 871.290 2.400 ;
        RECT 888.670 -4.800 889.230 2.400 ;
        RECT 906.610 -4.800 907.170 2.400 ;
        RECT 924.090 -4.800 924.650 2.400 ;
        RECT 942.030 -4.800 942.590 2.400 ;
        RECT 959.970 -4.800 960.530 2.400 ;
        RECT 977.910 -4.800 978.470 2.400 ;
        RECT 995.850 -4.800 996.410 2.400 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[0]
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 184.020 3466.000 187.020 3529.000 ;
        RECT 364.020 3466.000 367.020 3529.000 ;
        RECT 544.020 3466.000 547.020 3529.000 ;
        RECT 724.020 3466.000 727.020 3529.000 ;
        RECT 904.020 3466.000 907.020 3529.000 ;
        RECT 1084.020 3466.000 1087.020 3529.000 ;
        RECT 1264.020 3466.000 1267.020 3529.000 ;
        RECT 1444.020 3466.000 1447.020 3529.000 ;
        RECT 1624.020 3466.000 1627.020 3529.000 ;
        RECT 1804.020 3466.000 1807.020 3529.000 ;
        RECT 1984.020 3466.000 1987.020 3529.000 ;
        RECT 2164.020 3466.000 2167.020 3529.000 ;
        RECT 2344.020 3466.000 2347.020 3529.000 ;
        RECT 2524.020 3466.000 2527.020 3529.000 ;
        RECT 2704.020 3466.000 2707.020 3529.000 ;
        RECT 184.020 -9.320 187.020 54.000 ;
        RECT 364.020 -9.320 367.020 54.000 ;
        RECT 544.020 -9.320 547.020 54.000 ;
        RECT 724.020 -9.320 727.020 54.000 ;
        RECT 904.020 -9.320 907.020 54.000 ;
        RECT 1084.020 -9.320 1087.020 54.000 ;
        RECT 1264.020 -9.320 1267.020 54.000 ;
        RECT 1444.020 -9.320 1447.020 54.000 ;
        RECT 1624.020 -9.320 1627.020 54.000 ;
        RECT 1804.020 -9.320 1807.020 54.000 ;
        RECT 1984.020 -9.320 1987.020 54.000 ;
        RECT 2164.020 -9.320 2167.020 54.000 ;
        RECT 2344.020 -9.320 2347.020 54.000 ;
        RECT 2524.020 -9.320 2527.020 54.000 ;
        RECT 2704.020 -9.320 2707.020 54.000 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER M4M5_PR_C ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 54.000 3432.380 ;
        RECT 2866.000 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 54.000 3252.380 ;
        RECT 2866.000 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 54.000 3072.380 ;
        RECT 2866.000 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 54.000 2892.380 ;
        RECT 2866.000 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 54.000 2712.380 ;
        RECT 2866.000 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 54.000 2532.380 ;
        RECT 2866.000 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 54.000 2352.380 ;
        RECT 2866.000 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 54.000 2172.380 ;
        RECT 2866.000 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 54.000 1992.380 ;
        RECT 2866.000 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 54.000 1812.380 ;
        RECT 2866.000 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 54.000 1632.380 ;
        RECT 2866.000 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 54.000 1452.380 ;
        RECT 2866.000 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 54.000 1272.380 ;
        RECT 2866.000 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 54.000 1092.380 ;
        RECT 2866.000 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 54.000 912.380 ;
        RECT 2866.000 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 54.000 732.380 ;
        RECT 2866.000 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 54.000 552.380 ;
        RECT 2866.000 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 54.000 372.380 ;
        RECT 2866.000 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 54.000 192.380 ;
        RECT 2866.000 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 3466.000 97.020 3529.000 ;
        RECT 274.020 3466.000 277.020 3529.000 ;
        RECT 454.020 3466.000 457.020 3529.000 ;
        RECT 634.020 3466.000 637.020 3529.000 ;
        RECT 814.020 3466.000 817.020 3529.000 ;
        RECT 994.020 3466.000 997.020 3529.000 ;
        RECT 1174.020 3466.000 1177.020 3529.000 ;
        RECT 1354.020 3466.000 1357.020 3529.000 ;
        RECT 1534.020 3466.000 1537.020 3529.000 ;
        RECT 1714.020 3466.000 1717.020 3529.000 ;
        RECT 1894.020 3466.000 1897.020 3529.000 ;
        RECT 2074.020 3466.000 2077.020 3529.000 ;
        RECT 2254.020 3466.000 2257.020 3529.000 ;
        RECT 2434.020 3466.000 2437.020 3529.000 ;
        RECT 2614.020 3466.000 2617.020 3529.000 ;
        RECT 2794.020 3466.000 2797.020 3529.000 ;
        RECT 94.020 -9.320 97.020 54.000 ;
        RECT 274.020 -9.320 277.020 54.000 ;
        RECT 454.020 -9.320 457.020 54.000 ;
        RECT 634.020 -9.320 637.020 54.000 ;
        RECT 814.020 -9.320 817.020 54.000 ;
        RECT 994.020 -9.320 997.020 54.000 ;
        RECT 1174.020 -9.320 1177.020 54.000 ;
        RECT 1354.020 -9.320 1357.020 54.000 ;
        RECT 1534.020 -9.320 1537.020 54.000 ;
        RECT 1714.020 -9.320 1717.020 54.000 ;
        RECT 1894.020 -9.320 1897.020 54.000 ;
        RECT 2074.020 -9.320 2077.020 54.000 ;
        RECT 2254.020 -9.320 2257.020 54.000 ;
        RECT 2434.020 -9.320 2437.020 54.000 ;
        RECT 2614.020 -9.320 2617.020 54.000 ;
        RECT 2794.020 -9.320 2797.020 54.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER M4M5_PR_C ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 54.000 3342.380 ;
        RECT 2866.000 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 54.000 3162.380 ;
        RECT 2866.000 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 54.000 2982.380 ;
        RECT 2866.000 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 54.000 2802.380 ;
        RECT 2866.000 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 54.000 2622.380 ;
        RECT 2866.000 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 54.000 2442.380 ;
        RECT 2866.000 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 54.000 2262.380 ;
        RECT 2866.000 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 54.000 2082.380 ;
        RECT 2866.000 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 54.000 1902.380 ;
        RECT 2866.000 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 54.000 1722.380 ;
        RECT 2866.000 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 54.000 1542.380 ;
        RECT 2866.000 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 54.000 1362.380 ;
        RECT 2866.000 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 54.000 1182.380 ;
        RECT 2866.000 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 54.000 1002.380 ;
        RECT 2866.000 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 54.000 822.380 ;
        RECT 2866.000 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 54.000 642.380 ;
        RECT 2866.000 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 54.000 462.380 ;
        RECT 2866.000 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 54.000 282.380 ;
        RECT 2866.000 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 54.000 102.380 ;
        RECT 2866.000 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER M4M5_PR_C ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER M4M5_PR_C ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER M4M5_PR_C ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER M4M5_PR_C ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER M4M5_PR_C ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER M4M5_PR_C ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 95.825 331.675 2393.695 3466.000 ;
      LAYER met1 ;
        RECT 54.000 324.400 2866.000 3443.140 ;
      LAYER met2 ;
        RECT 54.840 54.000 2522.080 3466.000 ;
      LAYER met3 ;
        RECT 631.185 327.040 2414.935 2704.865 ;
      LAYER met4 ;
        RECT 94.020 54.000 2797.020 3466.000 ;
      LAYER met5 ;
        RECT 54.000 99.370 2866.000 3432.390 ;
  END
END user_project_wrapper
END LIBRARY

