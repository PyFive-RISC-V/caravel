VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 3005.380 BY 3594.740 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 66.810 2962.880 67.410 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 2412.810 2962.880 2413.410 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 2647.410 2962.880 2648.010 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 2882.010 2962.880 2882.610 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 3116.610 2962.880 3117.210 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 3351.210 2962.880 3351.810 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2922.110 3553.530 2922.390 3557.530 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2597.810 3553.530 2598.090 3557.530 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2273.510 3553.530 2273.790 3557.530 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1948.750 3553.530 1949.030 3557.530 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1624.450 3553.530 1624.730 3557.530 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 301.410 2962.880 302.010 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1300.150 3553.530 1300.430 3557.530 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 975.390 3553.530 975.670 3557.530 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 651.090 3553.530 651.370 3557.530 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 326.790 3553.530 327.070 3557.530 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 3520.530 46.880 3521.130 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 3232.890 46.880 3233.490 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 2945.930 46.880 2946.530 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 2658.290 46.880 2658.890 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 2371.330 46.880 2371.930 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 2083.690 46.880 2084.290 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 536.010 2962.880 536.610 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 1796.730 46.880 1797.330 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 770.610 2962.880 771.210 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 1005.210 2962.880 1005.810 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 1239.810 2962.880 1240.410 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 1474.410 2962.880 1475.010 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 1709.010 2962.880 1709.610 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 1943.610 2962.880 1944.210 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 2178.210 2962.880 2178.810 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 125.290 2962.880 125.890 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 2471.290 2962.880 2471.890 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 2707.020 2962.880 2707.170 ;
        RECT 2951.380 2706.720 2962.880 2707.020 ;
        RECT 2958.880 2706.570 2962.880 2706.720 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 2941.620 2962.880 2941.770 ;
        RECT 2951.380 2941.320 2962.880 2941.620 ;
        RECT 2958.880 2941.170 2962.880 2941.320 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 3176.220 2962.880 3176.370 ;
        RECT 2951.380 3175.920 2962.880 3176.220 ;
        RECT 2958.880 3175.770 2962.880 3175.920 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 3410.820 2962.880 3410.970 ;
        RECT 2951.380 3410.520 2962.880 3410.820 ;
        RECT 2958.880 3410.370 2962.880 3410.520 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2841.150 3553.530 2841.430 3557.530 ;
        RECT 2841.220 3540.740 2841.360 3553.530 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2516.850 3553.530 2517.130 3557.530 ;
        RECT 2516.920 3540.740 2517.060 3553.530 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2192.090 3553.530 2192.370 3557.530 ;
        RECT 2192.160 3540.740 2192.300 3553.530 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1867.790 3553.530 1868.070 3557.530 ;
        RECT 1867.860 3540.740 1868.000 3553.530 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1543.490 3553.530 1543.770 3557.530 ;
        RECT 1543.560 3540.740 1543.700 3553.530 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 359.890 2962.880 360.490 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1218.710 3542.490 1219.030 3542.550 ;
        RECT 2437.710 3542.490 2438.030 3542.550 ;
        RECT 1218.710 3542.350 2438.030 3542.490 ;
        RECT 1218.710 3542.290 1219.030 3542.350 ;
        RECT 2437.710 3542.290 2438.030 3542.350 ;
      LAYER via ;
        RECT 1218.740 3542.290 1219.000 3542.550 ;
        RECT 2437.740 3542.290 2438.000 3542.550 ;
      LAYER met2 ;
        RECT 1218.730 3553.530 1219.010 3557.530 ;
        RECT 1218.800 3542.580 1218.940 3553.530 ;
        RECT 1218.740 3542.260 1219.000 3542.580 ;
        RECT 2437.740 3542.260 2438.000 3542.580 ;
        RECT 2437.800 3540.740 2437.940 3542.260 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 894.410 3541.470 894.730 3541.530 ;
        RECT 2438.170 3541.470 2438.490 3541.530 ;
        RECT 894.410 3541.330 2438.490 3541.470 ;
        RECT 894.410 3541.270 894.730 3541.330 ;
        RECT 2438.170 3541.270 2438.490 3541.330 ;
      LAYER via ;
        RECT 894.440 3541.270 894.700 3541.530 ;
        RECT 2438.200 3541.270 2438.460 3541.530 ;
      LAYER met2 ;
        RECT 894.430 3553.530 894.710 3557.530 ;
        RECT 894.500 3541.560 894.640 3553.530 ;
        RECT 894.440 3541.240 894.700 3541.560 ;
        RECT 2438.200 3541.240 2438.460 3541.560 ;
        RECT 2438.260 3540.740 2438.400 3541.240 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 570.130 3553.530 570.410 3557.530 ;
        RECT 570.200 3540.740 570.340 3553.530 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 245.370 3553.530 245.650 3557.530 ;
        RECT 245.440 3540.740 245.580 3553.530 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 3448.900 46.880 3449.050 ;
        RECT 42.880 3448.600 54.000 3448.900 ;
        RECT 42.880 3448.450 46.880 3448.600 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 3161.940 46.880 3162.090 ;
        RECT 42.880 3161.640 54.000 3161.940 ;
        RECT 42.880 3161.490 46.880 3161.640 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 2874.300 46.880 2874.450 ;
        RECT 42.880 2874.000 54.000 2874.300 ;
        RECT 42.880 2873.850 46.880 2874.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 2586.890 46.880 2587.490 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 2299.250 46.880 2299.850 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 2012.290 46.880 2012.890 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 594.490 2962.880 595.090 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 1724.650 46.880 1725.250 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 1509.090 46.880 1509.690 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 1293.530 46.880 1294.130 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 1077.970 46.880 1078.570 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 862.410 46.880 863.010 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 647.530 46.880 648.130 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 431.970 46.880 432.570 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 42.880 216.410 46.880 217.010 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 829.090 2962.880 829.690 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 1063.690 2962.880 1064.290 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 1298.290 2962.880 1298.890 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 1532.890 2962.880 1533.490 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 1767.490 2962.880 1768.090 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 2002.090 2962.880 2002.690 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2958.880 2236.690 2962.880 2237.290 ;
    END
  END io_in[9]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2958.880 2823.980 2962.880 2824.130 ;
        RECT 2951.380 2823.680 2962.880 2823.980 ;
        RECT 2958.880 2823.530 2962.880 2823.680 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2958.880 3058.580 2962.880 3058.730 ;
        RECT 2951.380 3058.280 2962.880 3058.580 ;
        RECT 2958.880 3058.130 2962.880 3058.280 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2958.880 3293.180 2962.880 3293.330 ;
        RECT 2951.380 3292.880 2962.880 3293.180 ;
        RECT 2958.880 3292.730 2962.880 3292.880 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2958.880 3527.780 2962.880 3527.930 ;
        RECT 2951.380 3527.480 2962.880 3527.780 ;
        RECT 2958.880 3527.330 2962.880 3527.480 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2678.770 3553.530 2679.050 3557.530 ;
        RECT 2678.840 3540.740 2678.980 3553.530 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2354.470 3553.530 2354.750 3557.530 ;
        RECT 2354.540 3540.740 2354.680 3553.530 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.170 3553.530 2030.450 3557.530 ;
        RECT 2030.240 3540.740 2030.380 3553.530 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1705.410 3553.530 1705.690 3557.530 ;
        RECT 1705.480 3540.740 1705.620 3553.530 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1381.110 3553.530 1381.390 3557.530 ;
        RECT 1381.180 3540.740 1381.320 3553.530 ;
    END
  END io_oeb[19]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1056.790 3541.810 1057.110 3541.870 ;
        RECT 2431.270 3541.810 2431.590 3541.870 ;
        RECT 1056.790 3541.670 2431.590 3541.810 ;
        RECT 1056.790 3541.610 1057.110 3541.670 ;
        RECT 2431.270 3541.610 2431.590 3541.670 ;
      LAYER via ;
        RECT 1056.820 3541.610 1057.080 3541.870 ;
        RECT 2431.300 3541.610 2431.560 3541.870 ;
      LAYER met2 ;
        RECT 1056.810 3553.530 1057.090 3557.530 ;
        RECT 1056.880 3541.900 1057.020 3553.530 ;
        RECT 1056.820 3541.580 1057.080 3541.900 ;
        RECT 2431.300 3541.580 2431.560 3541.900 ;
        RECT 2431.360 3540.740 2431.500 3541.580 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 732.030 3540.790 732.350 3540.850 ;
        RECT 2433.110 3540.790 2433.430 3540.850 ;
        RECT 732.030 3540.740 2433.430 3540.790 ;
      LAYER via ;
        RECT 732.060 3540.740 732.320 3540.850 ;
        RECT 2433.140 3540.740 2433.400 3540.850 ;
      LAYER met2 ;
        RECT 732.050 3553.530 732.330 3557.530 ;
        RECT 732.120 3540.880 732.260 3553.530 ;
        RECT 732.060 3540.740 732.320 3540.880 ;
        RECT 2433.140 3540.740 2433.400 3540.880 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 407.750 3553.530 408.030 3557.530 ;
        RECT 407.820 3540.740 407.960 3553.530 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.450 3553.530 83.730 3557.530 ;
        RECT 83.520 3540.740 83.660 3553.530 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 42.880 3305.420 46.880 3305.570 ;
        RECT 42.880 3305.120 54.000 3305.420 ;
        RECT 42.880 3304.970 46.880 3305.120 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 42.880 3017.780 46.880 3017.930 ;
        RECT 42.880 3017.480 54.000 3017.780 ;
        RECT 42.880 3017.330 46.880 3017.480 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 42.880 2730.820 46.880 2730.970 ;
        RECT 42.880 2730.520 54.000 2730.820 ;
        RECT 42.880 2730.370 46.880 2730.520 ;
    END
  END io_oeb[26]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2958.880 2765.500 2962.880 2765.650 ;
        RECT 2951.380 2765.200 2962.880 2765.500 ;
        RECT 2958.880 2765.050 2962.880 2765.200 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2958.880 3000.100 2962.880 3000.250 ;
        RECT 2951.380 2999.800 2962.880 3000.100 ;
        RECT 2958.880 2999.650 2962.880 2999.800 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2958.880 3234.700 2962.880 3234.850 ;
        RECT 2951.380 3234.400 2962.880 3234.700 ;
        RECT 2958.880 3234.250 2962.880 3234.400 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2958.880 3469.300 2962.880 3469.450 ;
        RECT 2951.380 3469.000 2962.880 3469.300 ;
        RECT 2958.880 3468.850 2962.880 3469.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2760.190 3553.530 2760.470 3557.530 ;
        RECT 2760.260 3540.740 2760.400 3553.530 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2435.430 3553.530 2435.710 3557.530 ;
        RECT 2435.500 3542.660 2435.640 3553.530 ;
        RECT 2435.500 3542.520 2437.480 3542.660 ;
        RECT 2437.340 3540.740 2437.480 3542.520 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2111.130 3553.530 2111.410 3557.530 ;
        RECT 2111.200 3540.740 2111.340 3553.530 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1786.830 3553.530 1787.110 3557.530 ;
        RECT 1786.900 3540.740 1787.040 3553.530 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1462.070 3553.530 1462.350 3557.530 ;
        RECT 1462.140 3540.740 1462.280 3553.530 ;
    END
  END io_out[19]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1137.750 3542.150 1138.070 3542.210 ;
        RECT 2436.790 3542.150 2437.110 3542.210 ;
        RECT 1137.750 3542.010 2437.110 3542.150 ;
        RECT 1137.750 3541.950 1138.070 3542.010 ;
        RECT 2436.790 3541.950 2437.110 3542.010 ;
      LAYER via ;
        RECT 1137.780 3541.950 1138.040 3542.210 ;
        RECT 2436.820 3541.950 2437.080 3542.210 ;
      LAYER met2 ;
        RECT 1137.770 3553.530 1138.050 3557.530 ;
        RECT 1137.840 3542.240 1137.980 3553.530 ;
        RECT 1137.780 3541.920 1138.040 3542.240 ;
        RECT 2436.820 3541.920 2437.080 3542.240 ;
        RECT 2436.880 3540.740 2437.020 3541.920 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 813.450 3541.130 813.770 3541.190 ;
        RECT 2438.630 3541.130 2438.950 3541.190 ;
        RECT 813.450 3540.990 2438.950 3541.130 ;
        RECT 813.450 3540.930 813.770 3540.990 ;
        RECT 2438.630 3540.930 2438.950 3540.990 ;
      LAYER via ;
        RECT 813.480 3540.930 813.740 3541.190 ;
        RECT 2438.660 3540.930 2438.920 3541.190 ;
      LAYER met2 ;
        RECT 813.470 3553.530 813.750 3557.530 ;
        RECT 813.540 3541.220 813.680 3553.530 ;
        RECT 813.480 3540.900 813.740 3541.220 ;
        RECT 2438.660 3540.900 2438.920 3541.220 ;
        RECT 2438.720 3540.740 2438.860 3540.900 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 488.710 3553.530 488.990 3557.530 ;
        RECT 488.780 3540.740 488.920 3553.530 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 164.410 3553.530 164.690 3557.530 ;
        RECT 164.480 3540.740 164.620 3553.530 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 42.880 3377.500 46.880 3377.650 ;
        RECT 42.880 3377.200 54.000 3377.500 ;
        RECT 42.880 3377.050 46.880 3377.200 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 42.880 3089.860 46.880 3090.010 ;
        RECT 42.880 3089.560 54.000 3089.860 ;
        RECT 42.880 3089.410 46.880 3089.560 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 42.880 2802.900 46.880 2803.050 ;
        RECT 42.880 2802.600 54.000 2802.900 ;
        RECT 42.880 2802.450 46.880 2802.600 ;
    END
  END io_out[26]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 675.930 37.530 676.210 41.530 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2460.270 37.530 2460.550 41.530 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2477.750 37.530 2478.030 41.530 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2495.690 37.530 2495.970 41.530 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2513.630 37.530 2513.910 41.530 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2531.570 37.530 2531.850 41.530 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2549.050 37.530 2549.330 41.530 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2566.990 37.530 2567.270 41.530 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2584.930 37.530 2585.210 41.530 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2602.870 37.530 2603.150 41.530 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2620.810 37.530 2621.090 41.530 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 854.410 37.530 854.690 41.530 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2638.290 37.530 2638.570 41.530 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2656.230 37.530 2656.510 41.530 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2674.170 37.530 2674.450 41.530 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2692.110 37.530 2692.390 41.530 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2710.050 37.530 2710.330 41.530 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2727.530 37.530 2727.810 41.530 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2745.470 37.530 2745.750 41.530 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2763.410 37.530 2763.690 41.530 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2781.350 37.530 2781.630 41.530 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2798.830 37.530 2799.110 41.530 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 872.350 37.530 872.630 41.530 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2816.770 37.530 2817.050 41.530 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2834.710 37.530 2834.990 41.530 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2852.650 37.530 2852.930 41.530 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2870.590 37.530 2870.870 41.530 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2888.070 37.530 2888.350 41.530 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2906.010 37.530 2906.290 41.530 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2923.950 37.530 2924.230 41.530 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2941.890 37.530 2942.170 41.530 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 889.830 37.530 890.110 41.530 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 907.770 37.530 908.050 41.530 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 925.710 37.530 925.990 41.530 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 943.650 37.530 943.930 41.530 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 961.590 37.530 961.870 41.530 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 979.070 37.530 979.350 41.530 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 997.010 37.530 997.290 41.530 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1014.950 37.530 1015.230 41.530 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 693.870 37.530 694.150 41.530 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1032.890 37.530 1033.170 41.530 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1050.370 37.530 1050.650 41.530 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1068.310 37.530 1068.590 41.530 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1086.250 37.530 1086.530 41.530 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1104.190 37.530 1104.470 41.530 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1122.130 37.530 1122.410 41.530 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1139.610 37.530 1139.890 41.530 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1157.550 37.530 1157.830 41.530 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.490 37.530 1175.770 41.530 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1193.430 37.530 1193.710 41.530 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 711.810 37.530 712.090 41.530 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1211.370 37.530 1211.650 41.530 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1228.850 37.530 1229.130 41.530 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1246.790 37.530 1247.070 41.530 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1264.730 37.530 1265.010 41.530 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1282.670 37.530 1282.950 41.530 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1300.150 37.530 1300.430 41.530 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1318.090 37.530 1318.370 41.530 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1336.030 37.530 1336.310 41.530 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1353.970 37.530 1354.250 41.530 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1371.910 37.530 1372.190 41.530 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 729.290 37.530 729.570 41.530 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1389.390 37.530 1389.670 41.530 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1407.330 37.530 1407.610 41.530 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1425.270 37.530 1425.550 41.530 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1443.210 37.530 1443.490 41.530 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1461.150 37.530 1461.430 41.530 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1478.630 37.530 1478.910 41.530 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1496.570 37.530 1496.850 41.530 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1514.510 37.530 1514.790 41.530 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1532.450 37.530 1532.730 41.530 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1549.930 37.530 1550.210 41.530 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 747.230 37.530 747.510 41.530 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1567.870 37.530 1568.150 41.530 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1585.810 37.530 1586.090 41.530 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1603.750 37.530 1604.030 41.530 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1621.690 37.530 1621.970 41.530 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1639.170 37.530 1639.450 41.530 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1657.110 37.530 1657.390 41.530 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1675.050 37.530 1675.330 41.530 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1692.990 37.530 1693.270 41.530 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1710.930 37.530 1711.210 41.530 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1728.410 37.530 1728.690 41.530 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 765.170 37.530 765.450 41.530 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1746.350 37.530 1746.630 41.530 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1764.290 37.530 1764.570 41.530 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1782.230 37.530 1782.510 41.530 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1799.710 37.530 1799.990 41.530 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1817.650 37.530 1817.930 41.530 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1835.590 37.530 1835.870 41.530 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1853.530 37.530 1853.810 41.530 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1871.470 37.530 1871.750 41.530 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1888.950 37.530 1889.230 41.530 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1906.890 37.530 1907.170 41.530 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.110 37.530 783.390 41.530 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1924.830 37.530 1925.110 41.530 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1942.770 37.530 1943.050 41.530 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1960.710 37.530 1960.990 41.530 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1978.190 37.530 1978.470 41.530 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1996.130 37.530 1996.410 41.530 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2014.070 37.530 2014.350 41.530 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2032.010 37.530 2032.290 41.530 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2049.490 37.530 2049.770 41.530 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2067.430 37.530 2067.710 41.530 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2085.370 37.530 2085.650 41.530 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 800.590 37.530 800.870 41.530 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2103.310 37.530 2103.590 41.530 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2121.250 37.530 2121.530 41.530 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2138.730 37.530 2139.010 41.530 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2156.670 37.530 2156.950 41.530 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2174.610 37.530 2174.890 41.530 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2192.550 37.530 2192.830 41.530 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2210.490 37.530 2210.770 41.530 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2227.970 37.530 2228.250 41.530 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2245.910 37.530 2246.190 41.530 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2263.850 37.530 2264.130 41.530 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 818.530 37.530 818.810 41.530 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2281.790 37.530 2282.070 41.530 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2299.270 37.530 2299.550 41.530 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2317.210 37.530 2317.490 41.530 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2335.150 37.530 2335.430 41.530 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2353.090 37.530 2353.370 41.530 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2371.030 37.530 2371.310 41.530 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2388.510 37.530 2388.790 41.530 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2406.450 37.530 2406.730 41.530 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2424.390 37.530 2424.670 41.530 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2442.330 37.530 2442.610 41.530 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 836.470 37.530 836.750 41.530 ;
    END
  END la_data_in[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 687.890 37.530 688.170 41.530 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2471.770 37.530 2472.050 41.530 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2489.710 37.530 2489.990 41.530 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2507.650 37.530 2507.930 41.530 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2525.590 37.530 2525.870 41.530 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2543.530 37.530 2543.810 41.530 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2561.010 37.530 2561.290 41.530 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2578.950 37.530 2579.230 41.530 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2596.890 37.530 2597.170 41.530 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2614.830 37.530 2615.110 41.530 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2632.310 37.530 2632.590 41.530 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 866.370 37.530 866.650 41.530 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2650.250 37.530 2650.530 41.530 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2668.190 37.530 2668.470 41.530 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2686.130 37.530 2686.410 41.530 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2704.070 37.530 2704.350 41.530 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2721.550 37.530 2721.830 41.530 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2739.490 37.530 2739.770 41.530 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2757.430 37.530 2757.710 41.530 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2775.370 37.530 2775.650 41.530 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2793.310 37.530 2793.590 41.530 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2810.790 37.530 2811.070 41.530 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 883.850 37.530 884.130 41.530 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2828.730 37.530 2829.010 41.530 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2846.670 37.530 2846.950 41.530 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2864.610 37.530 2864.890 41.530 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2882.090 37.530 2882.370 41.530 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2900.030 37.530 2900.310 41.530 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2917.970 37.530 2918.250 41.530 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2935.910 37.530 2936.190 41.530 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2953.850 37.530 2954.130 41.530 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 901.790 37.530 902.070 41.530 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 919.730 37.530 920.010 41.530 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 937.670 37.530 937.950 41.530 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 955.610 37.530 955.890 41.530 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 973.090 37.530 973.370 41.530 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 991.030 37.530 991.310 41.530 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1008.970 37.530 1009.250 41.530 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1026.910 37.530 1027.190 41.530 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 705.830 37.530 706.110 41.530 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1044.850 37.530 1045.130 41.530 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1062.330 37.530 1062.610 41.530 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1080.270 37.530 1080.550 41.530 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1098.210 37.530 1098.490 41.530 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1116.150 37.530 1116.430 41.530 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1133.630 37.530 1133.910 41.530 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1151.570 37.530 1151.850 41.530 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1169.510 37.530 1169.790 41.530 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1187.450 37.530 1187.730 41.530 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1205.390 37.530 1205.670 41.530 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 723.310 37.530 723.590 41.530 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1222.870 37.530 1223.150 41.530 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1240.810 37.530 1241.090 41.530 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1258.750 37.530 1259.030 41.530 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1276.690 37.530 1276.970 41.530 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1294.630 37.530 1294.910 41.530 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1312.110 37.530 1312.390 41.530 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1330.050 37.530 1330.330 41.530 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1347.990 37.530 1348.270 41.530 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1365.930 37.530 1366.210 41.530 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1383.410 37.530 1383.690 41.530 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 741.250 37.530 741.530 41.530 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1401.350 37.530 1401.630 41.530 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1419.290 37.530 1419.570 41.530 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1437.230 37.530 1437.510 41.530 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1455.170 37.530 1455.450 41.530 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1472.650 37.530 1472.930 41.530 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1490.590 37.530 1490.870 41.530 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1508.530 37.530 1508.810 41.530 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1526.470 37.530 1526.750 41.530 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1544.410 37.530 1544.690 41.530 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1561.890 37.530 1562.170 41.530 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 759.190 37.530 759.470 41.530 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1579.830 37.530 1580.110 41.530 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1597.770 37.530 1598.050 41.530 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1615.710 37.530 1615.990 41.530 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1633.190 37.530 1633.470 41.530 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1651.130 37.530 1651.410 41.530 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1669.070 37.530 1669.350 41.530 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1687.010 37.530 1687.290 41.530 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1704.950 37.530 1705.230 41.530 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1722.430 37.530 1722.710 41.530 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1740.370 37.530 1740.650 41.530 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 777.130 37.530 777.410 41.530 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1758.310 37.530 1758.590 41.530 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1776.250 37.530 1776.530 41.530 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1794.190 37.530 1794.470 41.530 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1811.670 37.530 1811.950 41.530 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1829.610 37.530 1829.890 41.530 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1847.550 37.530 1847.830 41.530 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1865.490 37.530 1865.770 41.530 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1882.970 37.530 1883.250 41.530 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1900.910 37.530 1901.190 41.530 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1918.850 37.530 1919.130 41.530 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 795.070 37.530 795.350 41.530 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1936.790 37.530 1937.070 41.530 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1954.730 37.530 1955.010 41.530 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1972.210 37.530 1972.490 41.530 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1990.150 37.530 1990.430 41.530 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2008.090 37.530 2008.370 41.530 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2026.030 37.530 2026.310 41.530 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2043.970 37.530 2044.250 41.530 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2061.450 37.530 2061.730 41.530 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2079.390 37.530 2079.670 41.530 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2097.330 37.530 2097.610 41.530 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 812.550 37.530 812.830 41.530 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2115.270 37.530 2115.550 41.530 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2132.750 37.530 2133.030 41.530 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2150.690 37.530 2150.970 41.530 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2168.630 37.530 2168.910 41.530 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2186.570 37.530 2186.850 41.530 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2204.510 37.530 2204.790 41.530 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2221.990 37.530 2222.270 41.530 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2239.930 37.530 2240.210 41.530 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2257.870 37.530 2258.150 41.530 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2275.810 37.530 2276.090 41.530 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 830.490 37.530 830.770 41.530 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2293.750 37.530 2294.030 41.530 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2311.230 37.530 2311.510 41.530 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2329.170 37.530 2329.450 41.530 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2347.110 37.530 2347.390 41.530 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2365.050 37.530 2365.330 41.530 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2382.530 37.530 2382.810 41.530 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2400.470 37.530 2400.750 41.530 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2418.410 37.530 2418.690 41.530 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2436.350 37.530 2436.630 41.530 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2454.290 37.530 2454.570 41.530 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 848.430 37.530 848.710 41.530 ;
    END
  END la_oen[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2958.880 2589.380 2962.880 2589.530 ;
        RECT 2951.380 2589.080 2962.880 2589.380 ;
        RECT 2958.880 2588.930 2962.880 2589.080 ;
        RECT 2958.880 2530.900 2962.880 2531.050 ;
        RECT 2951.380 2530.600 2962.880 2530.900 ;
        RECT 2958.880 2530.450 2962.880 2530.600 ;
        RECT 42.880 2515.260 46.880 2515.410 ;
        RECT 42.880 2514.960 54.000 2515.260 ;
        RECT 42.880 2514.810 46.880 2514.960 ;
        RECT 42.880 2443.180 46.880 2443.330 ;
        RECT 42.880 2442.880 54.000 2443.180 ;
        RECT 42.880 2442.730 46.880 2442.880 ;
        RECT 2958.880 2354.780 2962.880 2354.930 ;
        RECT 2951.380 2354.480 2962.880 2354.780 ;
        RECT 2958.880 2354.330 2962.880 2354.480 ;
        RECT 2958.880 2296.300 2962.880 2296.450 ;
        RECT 2951.380 2296.000 2962.880 2296.300 ;
        RECT 2958.880 2295.850 2962.880 2296.000 ;
        RECT 42.880 2227.620 46.880 2227.770 ;
        RECT 42.880 2227.320 54.000 2227.620 ;
        RECT 42.880 2227.170 46.880 2227.320 ;
        RECT 42.880 2156.220 46.880 2156.370 ;
        RECT 42.880 2155.920 54.000 2156.220 ;
        RECT 42.880 2155.770 46.880 2155.920 ;
        RECT 2958.880 2120.180 2962.880 2120.330 ;
        RECT 2951.380 2119.880 2962.880 2120.180 ;
        RECT 2958.880 2119.730 2962.880 2119.880 ;
        RECT 2958.880 2061.700 2962.880 2061.850 ;
        RECT 2951.380 2061.400 2962.880 2061.700 ;
        RECT 2958.880 2061.250 2962.880 2061.400 ;
        RECT 42.880 1940.660 46.880 1940.810 ;
        RECT 42.880 1940.360 54.000 1940.660 ;
        RECT 42.880 1940.210 46.880 1940.360 ;
        RECT 2958.880 1885.580 2962.880 1885.730 ;
        RECT 2951.380 1885.280 2962.880 1885.580 ;
        RECT 2958.880 1885.130 2962.880 1885.280 ;
        RECT 42.880 1868.580 46.880 1868.730 ;
        RECT 42.880 1868.280 54.000 1868.580 ;
        RECT 42.880 1868.130 46.880 1868.280 ;
        RECT 2958.880 1827.100 2962.880 1827.250 ;
        RECT 2951.380 1826.800 2962.880 1827.100 ;
        RECT 2958.880 1826.650 2962.880 1826.800 ;
        RECT 42.880 1653.020 46.880 1653.170 ;
        RECT 42.880 1652.720 54.000 1653.020 ;
        RECT 42.880 1652.570 46.880 1652.720 ;
        RECT 2958.880 1650.980 2962.880 1651.130 ;
        RECT 2951.380 1650.680 2962.880 1650.980 ;
        RECT 2958.880 1650.530 2962.880 1650.680 ;
        RECT 2958.880 1591.820 2962.880 1591.970 ;
        RECT 2951.380 1591.520 2962.880 1591.820 ;
        RECT 2958.880 1591.370 2962.880 1591.520 ;
        RECT 42.880 1581.620 46.880 1581.770 ;
        RECT 42.880 1581.320 54.000 1581.620 ;
        RECT 42.880 1581.170 46.880 1581.320 ;
        RECT 42.880 1438.140 46.880 1438.290 ;
        RECT 42.880 1437.840 54.000 1438.140 ;
        RECT 42.880 1437.690 46.880 1437.840 ;
        RECT 2958.880 1416.380 2962.880 1416.530 ;
        RECT 2951.380 1416.080 2962.880 1416.380 ;
        RECT 2958.880 1415.930 2962.880 1416.080 ;
        RECT 42.880 1366.060 46.880 1366.210 ;
        RECT 42.880 1365.760 54.000 1366.060 ;
        RECT 42.880 1365.610 46.880 1365.760 ;
        RECT 2958.880 1357.220 2962.880 1357.370 ;
        RECT 2951.380 1356.920 2962.880 1357.220 ;
        RECT 2958.880 1356.770 2962.880 1356.920 ;
        RECT 42.880 1222.580 46.880 1222.730 ;
        RECT 42.880 1222.280 54.000 1222.580 ;
        RECT 42.880 1222.130 46.880 1222.280 ;
        RECT 2958.880 1181.780 2962.880 1181.930 ;
        RECT 2951.380 1181.480 2962.880 1181.780 ;
        RECT 2958.880 1181.330 2962.880 1181.480 ;
        RECT 42.880 1150.500 46.880 1150.650 ;
        RECT 42.880 1150.200 54.000 1150.500 ;
        RECT 42.880 1150.050 46.880 1150.200 ;
        RECT 2958.880 1122.620 2962.880 1122.770 ;
        RECT 2951.380 1122.320 2962.880 1122.620 ;
        RECT 2958.880 1122.170 2962.880 1122.320 ;
        RECT 42.880 1007.020 46.880 1007.170 ;
        RECT 42.880 1006.720 54.000 1007.020 ;
        RECT 42.880 1006.570 46.880 1006.720 ;
        RECT 2958.880 947.180 2962.880 947.330 ;
        RECT 2951.380 946.880 2962.880 947.180 ;
        RECT 2958.880 946.730 2962.880 946.880 ;
        RECT 42.880 934.940 46.880 935.090 ;
        RECT 42.880 934.640 54.000 934.940 ;
        RECT 42.880 934.490 46.880 934.640 ;
        RECT 2958.880 888.020 2962.880 888.170 ;
        RECT 2951.380 887.720 2962.880 888.020 ;
        RECT 2958.880 887.570 2962.880 887.720 ;
        RECT 42.880 791.460 46.880 791.610 ;
        RECT 42.880 791.160 54.000 791.460 ;
        RECT 42.880 791.010 46.880 791.160 ;
        RECT 42.880 719.380 46.880 719.530 ;
        RECT 42.880 719.080 54.000 719.380 ;
        RECT 42.880 718.930 46.880 719.080 ;
        RECT 2958.880 711.900 2962.880 712.050 ;
        RECT 2951.380 711.600 2962.880 711.900 ;
        RECT 2958.880 711.450 2962.880 711.600 ;
        RECT 2958.880 653.420 2962.880 653.570 ;
        RECT 2951.380 653.120 2962.880 653.420 ;
        RECT 2958.880 652.970 2962.880 653.120 ;
        RECT 42.880 575.900 46.880 576.050 ;
        RECT 42.880 575.600 54.000 575.900 ;
        RECT 42.880 575.450 46.880 575.600 ;
        RECT 42.880 503.820 46.880 503.970 ;
        RECT 42.880 503.520 54.000 503.820 ;
        RECT 42.880 503.370 46.880 503.520 ;
        RECT 2958.880 477.300 2962.880 477.450 ;
        RECT 2951.380 477.000 2962.880 477.300 ;
        RECT 2958.880 476.850 2962.880 477.000 ;
        RECT 2958.880 418.820 2962.880 418.970 ;
        RECT 2951.380 418.520 2962.880 418.820 ;
        RECT 2958.880 418.370 2962.880 418.520 ;
        RECT 42.880 360.340 46.880 360.490 ;
        RECT 42.880 360.040 54.000 360.340 ;
        RECT 42.880 359.890 46.880 360.040 ;
        RECT 42.880 288.260 46.880 288.410 ;
        RECT 42.880 287.960 54.000 288.260 ;
        RECT 42.880 287.810 46.880 287.960 ;
        RECT 2958.880 242.700 2962.880 242.850 ;
        RECT 2951.380 242.400 2962.880 242.700 ;
        RECT 2958.880 242.250 2962.880 242.400 ;
        RECT 2958.880 184.220 2962.880 184.370 ;
        RECT 2951.380 183.920 2962.880 184.220 ;
        RECT 2958.880 183.770 2962.880 183.920 ;
        RECT 42.880 144.780 46.880 144.930 ;
        RECT 42.880 144.480 54.000 144.780 ;
        RECT 42.880 144.330 46.880 144.480 ;
        RECT 42.880 73.380 46.880 73.530 ;
        RECT 42.880 73.080 54.000 73.380 ;
        RECT 42.880 72.930 46.880 73.080 ;
    END
  END io_oeb[0]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2959.830 37.530 2960.110 41.530 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 49.390 362.130 49.710 362.190 ;
        RECT 49.390 361.990 54.000 362.130 ;
        RECT 49.390 361.930 49.710 361.990 ;
        RECT 45.710 54.090 46.030 54.150 ;
        RECT 49.390 54.090 49.710 54.150 ;
        RECT 45.710 53.950 49.710 54.090 ;
        RECT 45.710 53.890 46.030 53.950 ;
        RECT 49.390 53.890 49.710 53.950 ;
      LAYER via ;
        RECT 49.420 361.930 49.680 362.190 ;
        RECT 45.740 53.890 46.000 54.150 ;
        RECT 49.420 53.890 49.680 54.150 ;
      LAYER met2 ;
        RECT 49.420 361.900 49.680 362.220 ;
        RECT 49.480 54.180 49.620 361.900 ;
        RECT 45.740 53.860 46.000 54.180 ;
        RECT 49.420 53.860 49.680 54.180 ;
        RECT 45.800 41.530 45.940 53.860 ;
        RECT 45.730 37.530 46.010 41.530 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 51.230 54.770 51.550 54.830 ;
        RECT 51.230 54.630 54.000 54.770 ;
        RECT 51.230 54.570 51.550 54.630 ;
      LAYER via ;
        RECT 51.260 54.570 51.520 54.830 ;
      LAYER met2 ;
        RECT 51.260 54.540 51.520 54.860 ;
        RECT 51.320 41.530 51.460 54.540 ;
        RECT 51.250 37.530 51.530 41.530 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 57.300 41.530 57.440 54.000 ;
        RECT 57.230 37.530 57.510 41.530 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.220 41.530 81.360 54.000 ;
        RECT 81.150 37.530 81.430 41.530 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 283.620 41.530 283.760 54.000 ;
        RECT 283.550 37.530 283.830 41.530 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 301.100 41.530 301.240 54.000 ;
        RECT 301.030 37.530 301.310 41.530 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.040 41.530 319.180 54.000 ;
        RECT 318.970 37.530 319.250 41.530 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 336.980 41.530 337.120 54.000 ;
        RECT 336.910 37.530 337.190 41.530 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 354.920 41.530 355.060 54.000 ;
        RECT 354.850 37.530 355.130 41.530 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 372.860 41.530 373.000 54.000 ;
        RECT 372.790 37.530 373.070 41.530 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.340 41.530 390.480 54.000 ;
        RECT 390.270 37.530 390.550 41.530 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 408.280 41.530 408.420 54.000 ;
        RECT 408.210 37.530 408.490 41.530 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 426.220 41.530 426.360 54.000 ;
        RECT 426.150 37.530 426.430 41.530 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 444.160 41.530 444.300 54.000 ;
        RECT 444.090 37.530 444.370 41.530 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.140 41.530 105.280 54.000 ;
        RECT 105.070 37.530 105.350 41.530 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 462.100 41.530 462.240 54.000 ;
        RECT 462.030 37.530 462.310 41.530 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 479.580 41.530 479.720 54.000 ;
        RECT 479.510 37.530 479.790 41.530 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 497.520 41.530 497.660 54.000 ;
        RECT 497.450 37.530 497.730 41.530 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 515.370 53.070 515.690 53.130 ;
        RECT 518.590 53.070 518.910 53.130 ;
        RECT 515.370 52.930 518.910 53.070 ;
        RECT 515.370 52.870 515.690 52.930 ;
        RECT 518.590 52.870 518.910 52.930 ;
      LAYER via ;
        RECT 515.400 52.870 515.660 53.130 ;
        RECT 518.620 52.870 518.880 53.130 ;
      LAYER met2 ;
        RECT 518.680 53.160 518.820 54.000 ;
        RECT 515.400 52.840 515.660 53.160 ;
        RECT 518.620 52.840 518.880 53.160 ;
        RECT 515.460 41.530 515.600 52.840 ;
        RECT 515.390 37.530 515.670 41.530 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 533.400 41.530 533.540 54.000 ;
        RECT 533.330 37.530 533.610 41.530 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 550.880 41.530 551.020 54.000 ;
        RECT 550.810 37.530 551.090 41.530 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 568.820 41.530 568.960 54.000 ;
        RECT 568.750 37.530 569.030 41.530 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 586.760 41.530 586.900 54.000 ;
        RECT 586.690 37.530 586.970 41.530 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 604.700 41.530 604.840 54.000 ;
        RECT 604.630 37.530 604.910 41.530 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 622.640 41.530 622.780 54.000 ;
        RECT 622.570 37.530 622.850 41.530 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.060 41.530 129.200 54.000 ;
        RECT 128.990 37.530 129.270 41.530 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 640.030 52.730 640.350 52.790 ;
        RECT 642.790 52.730 643.110 52.790 ;
        RECT 640.030 52.590 643.110 52.730 ;
        RECT 640.030 52.530 640.350 52.590 ;
        RECT 642.790 52.530 643.110 52.590 ;
      LAYER via ;
        RECT 640.060 52.530 640.320 52.790 ;
        RECT 642.820 52.530 643.080 52.790 ;
      LAYER met2 ;
        RECT 642.880 52.820 643.020 54.000 ;
        RECT 640.060 52.500 640.320 52.820 ;
        RECT 642.820 52.500 643.080 52.820 ;
        RECT 640.120 41.530 640.260 52.500 ;
        RECT 640.050 37.530 640.330 41.530 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 658.060 41.530 658.200 54.000 ;
        RECT 657.990 37.530 658.270 41.530 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 152.520 41.530 152.660 54.000 ;
        RECT 152.450 37.530 152.730 41.530 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.440 41.530 176.580 54.000 ;
        RECT 176.370 37.530 176.650 41.530 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 194.380 41.530 194.520 54.000 ;
        RECT 194.310 37.530 194.590 41.530 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 212.320 41.530 212.460 54.000 ;
        RECT 212.250 37.530 212.530 41.530 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 229.800 41.530 229.940 54.000 ;
        RECT 229.730 37.530 230.010 41.530 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 247.740 41.530 247.880 54.000 ;
        RECT 247.670 37.530 247.950 41.530 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 265.680 41.530 265.820 54.000 ;
        RECT 265.610 37.530 265.890 41.530 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.280 41.530 63.420 54.000 ;
        RECT 63.210 37.530 63.490 41.530 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 87.110 53.950 91.110 54.000 ;
        RECT 87.110 53.890 87.430 53.950 ;
        RECT 90.790 53.890 91.110 53.950 ;
      LAYER via ;
        RECT 87.140 53.890 87.400 54.000 ;
        RECT 90.820 53.890 91.080 54.000 ;
      LAYER met2 ;
        RECT 87.140 53.860 87.400 54.000 ;
        RECT 90.820 53.860 91.080 54.000 ;
        RECT 87.200 41.530 87.340 53.860 ;
        RECT 87.130 37.530 87.410 41.530 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 289.600 41.530 289.740 54.000 ;
        RECT 289.530 37.530 289.810 41.530 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 307.080 41.530 307.220 54.000 ;
        RECT 307.010 37.530 307.290 41.530 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 325.020 41.530 325.160 54.000 ;
        RECT 324.950 37.530 325.230 41.530 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 342.960 41.530 343.100 54.000 ;
        RECT 342.890 37.530 343.170 41.530 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 360.900 41.530 361.040 54.000 ;
        RECT 360.830 37.530 361.110 41.530 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 378.840 41.530 378.980 54.000 ;
        RECT 378.770 37.530 379.050 41.530 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 396.320 41.530 396.460 54.000 ;
        RECT 396.250 37.530 396.530 41.530 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 414.260 41.530 414.400 54.000 ;
        RECT 414.190 37.530 414.470 41.530 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 432.110 53.950 436.110 54.000 ;
        RECT 432.110 53.890 432.430 53.950 ;
        RECT 435.790 53.890 436.110 53.950 ;
      LAYER via ;
        RECT 432.140 53.890 432.400 54.000 ;
        RECT 435.820 53.890 436.080 54.000 ;
      LAYER met2 ;
        RECT 432.140 53.860 432.400 54.000 ;
        RECT 435.820 53.860 436.080 54.000 ;
        RECT 432.200 41.530 432.340 53.860 ;
        RECT 432.130 37.530 432.410 41.530 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 450.140 41.530 450.280 54.000 ;
        RECT 450.070 37.530 450.350 41.530 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.120 41.530 111.260 54.000 ;
        RECT 111.050 37.530 111.330 41.530 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 467.620 41.530 467.760 54.000 ;
        RECT 467.550 37.530 467.830 41.530 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 485.560 41.530 485.700 54.000 ;
        RECT 485.490 37.530 485.770 41.530 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 503.500 41.530 503.640 54.000 ;
        RECT 503.430 37.530 503.710 41.530 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 521.440 41.530 521.580 54.000 ;
        RECT 521.370 37.530 521.650 41.530 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 539.380 41.530 539.520 54.000 ;
        RECT 539.310 37.530 539.590 41.530 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 556.860 41.530 557.000 54.000 ;
        RECT 556.790 37.530 557.070 41.530 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 574.800 41.530 574.940 54.000 ;
        RECT 574.730 37.530 575.010 41.530 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 592.740 41.530 592.880 54.000 ;
        RECT 592.670 37.530 592.950 41.530 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 610.680 41.530 610.820 54.000 ;
        RECT 610.610 37.530 610.890 41.530 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 628.620 41.530 628.760 54.000 ;
        RECT 628.550 37.530 628.830 41.530 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.580 41.530 134.720 54.000 ;
        RECT 134.510 37.530 134.790 41.530 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 646.100 41.530 646.240 54.000 ;
        RECT 646.030 37.530 646.310 41.530 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 664.040 41.530 664.180 54.000 ;
        RECT 663.970 37.530 664.250 41.530 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 158.500 41.530 158.640 54.000 ;
        RECT 158.430 37.530 158.710 41.530 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 182.420 41.530 182.560 54.000 ;
        RECT 182.350 37.530 182.630 41.530 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 200.360 41.530 200.500 54.000 ;
        RECT 200.290 37.530 200.570 41.530 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.840 41.530 217.980 54.000 ;
        RECT 217.770 37.530 218.050 41.530 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 235.780 41.530 235.920 54.000 ;
        RECT 235.710 37.530 235.990 41.530 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 253.720 41.530 253.860 54.000 ;
        RECT 253.650 37.530 253.930 41.530 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 271.660 41.530 271.800 54.000 ;
        RECT 271.590 37.530 271.870 41.530 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.180 41.530 93.320 54.000 ;
        RECT 93.110 37.530 93.390 41.530 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 295.580 41.530 295.720 54.000 ;
        RECT 295.510 37.530 295.790 41.530 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 313.060 41.530 313.200 54.000 ;
        RECT 312.990 37.530 313.270 41.530 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 331.000 41.530 331.140 54.000 ;
        RECT 330.930 37.530 331.210 41.530 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 348.940 41.530 349.080 54.000 ;
        RECT 348.870 37.530 349.150 41.530 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 366.880 41.530 367.020 54.000 ;
        RECT 366.810 37.530 367.090 41.530 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 384.360 41.530 384.500 54.000 ;
        RECT 384.290 37.530 384.570 41.530 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 402.300 41.530 402.440 54.000 ;
        RECT 402.230 37.530 402.510 41.530 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 420.240 41.530 420.380 54.000 ;
        RECT 420.170 37.530 420.450 41.530 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 438.180 41.530 438.320 54.000 ;
        RECT 438.110 37.530 438.390 41.530 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 456.120 41.530 456.260 54.000 ;
        RECT 456.050 37.530 456.330 41.530 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.100 41.530 117.240 54.000 ;
        RECT 117.030 37.530 117.310 41.530 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 473.510 53.950 477.510 54.000 ;
        RECT 473.510 53.890 473.830 53.950 ;
        RECT 477.190 53.890 477.510 53.950 ;
      LAYER via ;
        RECT 473.540 53.890 473.800 54.000 ;
        RECT 477.220 53.890 477.480 54.000 ;
      LAYER met2 ;
        RECT 473.540 53.860 473.800 54.000 ;
        RECT 477.220 53.860 477.480 54.000 ;
        RECT 473.600 41.530 473.740 53.860 ;
        RECT 473.530 37.530 473.810 41.530 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 491.540 41.530 491.680 54.000 ;
        RECT 491.470 37.530 491.750 41.530 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 509.480 41.530 509.620 54.000 ;
        RECT 509.410 37.530 509.690 41.530 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 527.420 41.530 527.560 54.000 ;
        RECT 527.350 37.530 527.630 41.530 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 545.360 41.530 545.500 54.000 ;
        RECT 545.290 37.530 545.570 41.530 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 562.840 41.530 562.980 54.000 ;
        RECT 562.770 37.530 563.050 41.530 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 580.780 41.530 580.920 54.000 ;
        RECT 580.710 37.530 580.990 41.530 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 598.720 41.530 598.860 54.000 ;
        RECT 598.650 37.530 598.930 41.530 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 616.660 41.530 616.800 54.000 ;
        RECT 616.590 37.530 616.870 41.530 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 634.140 41.530 634.280 54.000 ;
        RECT 634.070 37.530 634.350 41.530 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 140.560 41.530 140.700 54.000 ;
        RECT 140.490 37.530 140.770 41.530 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 652.080 41.530 652.220 54.000 ;
        RECT 652.010 37.530 652.290 41.530 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 670.480 42.020 670.620 54.000 ;
        RECT 670.020 41.880 670.620 42.020 ;
        RECT 670.020 41.530 670.160 41.880 ;
        RECT 669.950 37.530 670.230 41.530 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 164.480 41.530 164.620 54.000 ;
        RECT 164.410 37.530 164.690 41.530 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 188.400 41.530 188.540 54.000 ;
        RECT 188.330 37.530 188.610 41.530 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 206.340 41.530 206.480 54.000 ;
        RECT 206.270 37.530 206.550 41.530 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 223.820 41.530 223.960 54.000 ;
        RECT 223.750 37.530 224.030 41.530 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 241.760 41.530 241.900 54.000 ;
        RECT 241.690 37.530 241.970 41.530 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 259.700 41.530 259.840 54.000 ;
        RECT 259.630 37.530 259.910 41.530 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 277.640 41.530 277.780 54.000 ;
        RECT 277.570 37.530 277.850 41.530 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.160 41.530 99.300 54.000 ;
        RECT 99.090 37.530 99.370 41.530 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.080 41.530 123.220 54.000 ;
        RECT 123.010 37.530 123.290 41.530 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 146.540 41.530 146.680 54.000 ;
        RECT 146.470 37.530 146.750 41.530 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.460 41.530 170.600 54.000 ;
        RECT 170.390 37.530 170.670 41.530 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.180 42.020 70.320 54.000 ;
        RECT 69.260 41.880 70.320 42.020 ;
        RECT 69.260 41.530 69.400 41.880 ;
        RECT 69.190 37.530 69.470 41.530 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.080 42.020 77.220 54.000 ;
        RECT 75.240 41.880 77.220 42.020 ;
        RECT 75.240 41.530 75.380 41.880 ;
        RECT 75.170 37.530 75.450 41.530 ;
    END
  END wbs_we_i
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 681.890 51.710 682.210 51.770 ;
        RECT 696.610 51.710 696.930 51.770 ;
        RECT 699.830 51.710 700.150 51.770 ;
        RECT 717.310 51.710 717.630 51.770 ;
        RECT 735.250 51.710 735.570 51.770 ;
        RECT 753.190 51.710 753.510 51.770 ;
        RECT 771.130 51.710 771.450 51.770 ;
        RECT 789.070 51.710 789.390 51.770 ;
        RECT 806.550 51.710 806.870 51.770 ;
        RECT 824.490 51.710 824.810 51.770 ;
        RECT 842.430 51.710 842.750 51.770 ;
        RECT 860.370 51.710 860.690 51.770 ;
        RECT 878.310 51.710 878.630 51.770 ;
        RECT 895.790 51.710 896.110 51.770 ;
        RECT 913.730 51.710 914.050 51.770 ;
        RECT 931.670 51.710 931.990 51.770 ;
        RECT 949.610 51.710 949.930 51.770 ;
        RECT 967.090 51.710 967.410 51.770 ;
        RECT 985.030 51.710 985.350 51.770 ;
        RECT 1002.970 51.710 1003.290 51.770 ;
        RECT 1020.910 51.710 1021.230 51.770 ;
        RECT 1038.850 51.710 1039.170 51.770 ;
        RECT 1056.330 51.710 1056.650 51.770 ;
        RECT 1074.270 51.710 1074.590 51.770 ;
        RECT 1092.210 51.710 1092.530 51.770 ;
        RECT 1110.150 51.710 1110.470 51.770 ;
        RECT 1128.090 51.710 1128.410 51.770 ;
        RECT 1145.570 51.710 1145.890 51.770 ;
        RECT 1163.510 51.710 1163.830 51.770 ;
        RECT 1181.450 51.710 1181.770 51.770 ;
        RECT 1199.390 51.710 1199.710 51.770 ;
        RECT 1216.870 51.710 1217.190 51.770 ;
        RECT 1234.810 51.710 1235.130 51.770 ;
        RECT 1252.750 51.710 1253.070 51.770 ;
        RECT 1270.690 51.710 1271.010 51.770 ;
        RECT 1288.630 51.710 1288.950 51.770 ;
        RECT 1306.110 51.710 1306.430 51.770 ;
        RECT 1324.050 51.710 1324.370 51.770 ;
        RECT 1341.990 51.710 1342.310 51.770 ;
        RECT 1359.930 51.710 1360.250 51.770 ;
        RECT 1377.870 51.710 1378.190 51.770 ;
        RECT 1395.350 51.710 1395.670 51.770 ;
        RECT 1413.290 51.710 1413.610 51.770 ;
        RECT 1431.230 51.710 1431.550 51.770 ;
        RECT 1449.170 51.710 1449.490 51.770 ;
        RECT 1466.650 51.710 1466.970 51.770 ;
        RECT 1484.590 51.710 1484.910 51.770 ;
        RECT 1502.530 51.710 1502.850 51.770 ;
        RECT 1520.470 51.710 1520.790 51.770 ;
        RECT 1538.410 51.710 1538.730 51.770 ;
        RECT 1555.890 51.710 1556.210 51.770 ;
        RECT 1573.830 51.710 1574.150 51.770 ;
        RECT 1591.770 51.710 1592.090 51.770 ;
        RECT 1609.710 51.710 1610.030 51.770 ;
        RECT 1627.650 51.710 1627.970 51.770 ;
        RECT 1645.130 51.710 1645.450 51.770 ;
        RECT 1663.070 51.710 1663.390 51.770 ;
        RECT 1681.010 51.710 1681.330 51.770 ;
        RECT 1698.950 51.710 1699.270 51.770 ;
        RECT 1716.430 51.710 1716.750 51.770 ;
        RECT 1734.370 51.710 1734.690 51.770 ;
        RECT 1752.310 51.710 1752.630 51.770 ;
        RECT 1770.250 51.710 1770.570 51.770 ;
        RECT 1788.190 51.710 1788.510 51.770 ;
        RECT 1805.670 51.710 1805.990 51.770 ;
        RECT 1823.610 51.710 1823.930 51.770 ;
        RECT 1841.550 51.710 1841.870 51.770 ;
        RECT 1859.490 51.710 1859.810 51.770 ;
        RECT 1877.430 51.710 1877.750 51.770 ;
        RECT 1894.910 51.710 1895.230 51.770 ;
        RECT 1912.850 51.710 1913.170 51.770 ;
        RECT 1930.790 51.710 1931.110 51.770 ;
        RECT 1948.730 51.710 1949.050 51.770 ;
        RECT 1966.210 51.710 1966.530 51.770 ;
        RECT 1984.150 51.710 1984.470 51.770 ;
        RECT 2002.090 51.710 2002.410 51.770 ;
        RECT 2020.030 51.710 2020.350 51.770 ;
        RECT 2037.970 51.710 2038.290 51.770 ;
        RECT 2055.450 51.710 2055.770 51.770 ;
        RECT 2073.390 51.710 2073.710 51.770 ;
        RECT 2091.330 51.710 2091.650 51.770 ;
        RECT 2109.270 51.710 2109.590 51.770 ;
        RECT 2127.210 51.710 2127.530 51.770 ;
        RECT 2144.690 51.710 2145.010 51.770 ;
        RECT 2162.630 51.710 2162.950 51.770 ;
        RECT 2180.570 51.710 2180.890 51.770 ;
        RECT 2198.510 51.710 2198.830 51.770 ;
        RECT 2215.990 51.710 2216.310 51.770 ;
        RECT 2233.930 51.710 2234.250 51.770 ;
        RECT 2251.870 51.710 2252.190 51.770 ;
        RECT 2269.810 51.710 2270.130 51.770 ;
        RECT 2287.750 51.710 2288.070 51.770 ;
        RECT 2305.230 51.710 2305.550 51.770 ;
        RECT 2323.170 51.710 2323.490 51.770 ;
        RECT 2341.110 51.710 2341.430 51.770 ;
        RECT 2359.050 51.710 2359.370 51.770 ;
        RECT 2376.990 51.710 2377.310 51.770 ;
        RECT 2394.470 51.710 2394.790 51.770 ;
        RECT 2412.410 51.710 2412.730 51.770 ;
        RECT 2430.350 51.710 2430.670 51.770 ;
        RECT 2448.290 51.710 2448.610 51.770 ;
        RECT 2465.770 51.710 2466.090 51.770 ;
        RECT 2483.710 51.710 2484.030 51.770 ;
        RECT 2501.650 51.710 2501.970 51.770 ;
        RECT 2519.590 51.710 2519.910 51.770 ;
        RECT 2537.530 51.710 2537.850 51.770 ;
        RECT 2555.010 51.710 2555.330 51.770 ;
        RECT 2572.950 51.710 2573.270 51.770 ;
        RECT 2590.890 51.710 2591.210 51.770 ;
        RECT 2608.830 51.710 2609.150 51.770 ;
        RECT 2626.770 51.710 2627.090 51.770 ;
        RECT 2644.250 51.710 2644.570 51.770 ;
        RECT 2662.190 51.710 2662.510 51.770 ;
        RECT 2680.130 51.710 2680.450 51.770 ;
        RECT 2698.070 51.710 2698.390 51.770 ;
        RECT 2715.550 51.710 2715.870 51.770 ;
        RECT 2733.490 51.710 2733.810 51.770 ;
        RECT 2751.430 51.710 2751.750 51.770 ;
        RECT 2769.370 51.710 2769.690 51.770 ;
        RECT 2787.310 51.710 2787.630 51.770 ;
        RECT 2804.790 51.710 2805.110 51.770 ;
        RECT 2822.730 51.710 2823.050 51.770 ;
        RECT 2840.670 51.710 2840.990 51.770 ;
        RECT 2858.610 51.710 2858.930 51.770 ;
        RECT 2876.550 51.710 2876.870 51.770 ;
        RECT 2894.030 51.710 2894.350 51.770 ;
        RECT 2911.970 51.710 2912.290 51.770 ;
        RECT 2929.910 51.710 2930.230 51.770 ;
        RECT 2947.850 51.710 2948.170 51.770 ;
        RECT 681.890 51.570 2948.170 51.710 ;
        RECT 681.890 51.510 682.210 51.570 ;
        RECT 696.610 51.510 696.930 51.570 ;
        RECT 699.830 51.510 700.150 51.570 ;
        RECT 717.310 51.510 717.630 51.570 ;
        RECT 735.250 51.510 735.570 51.570 ;
        RECT 753.190 51.510 753.510 51.570 ;
        RECT 771.130 51.510 771.450 51.570 ;
        RECT 789.070 51.510 789.390 51.570 ;
        RECT 806.550 51.510 806.870 51.570 ;
        RECT 824.490 51.510 824.810 51.570 ;
        RECT 842.430 51.510 842.750 51.570 ;
        RECT 860.370 51.510 860.690 51.570 ;
        RECT 878.310 51.510 878.630 51.570 ;
        RECT 895.790 51.510 896.110 51.570 ;
        RECT 913.730 51.510 914.050 51.570 ;
        RECT 931.670 51.510 931.990 51.570 ;
        RECT 949.610 51.510 949.930 51.570 ;
        RECT 967.090 51.510 967.410 51.570 ;
        RECT 985.030 51.510 985.350 51.570 ;
        RECT 1002.970 51.510 1003.290 51.570 ;
        RECT 1020.910 51.510 1021.230 51.570 ;
        RECT 1038.850 51.510 1039.170 51.570 ;
        RECT 1056.330 51.510 1056.650 51.570 ;
        RECT 1074.270 51.510 1074.590 51.570 ;
        RECT 1092.210 51.510 1092.530 51.570 ;
        RECT 1110.150 51.510 1110.470 51.570 ;
        RECT 1128.090 51.510 1128.410 51.570 ;
        RECT 1145.570 51.510 1145.890 51.570 ;
        RECT 1163.510 51.510 1163.830 51.570 ;
        RECT 1181.450 51.510 1181.770 51.570 ;
        RECT 1199.390 51.510 1199.710 51.570 ;
        RECT 1216.870 51.510 1217.190 51.570 ;
        RECT 1234.810 51.510 1235.130 51.570 ;
        RECT 1252.750 51.510 1253.070 51.570 ;
        RECT 1270.690 51.510 1271.010 51.570 ;
        RECT 1288.630 51.510 1288.950 51.570 ;
        RECT 1306.110 51.510 1306.430 51.570 ;
        RECT 1324.050 51.510 1324.370 51.570 ;
        RECT 1341.990 51.510 1342.310 51.570 ;
        RECT 1359.930 51.510 1360.250 51.570 ;
        RECT 1377.870 51.510 1378.190 51.570 ;
        RECT 1395.350 51.510 1395.670 51.570 ;
        RECT 1413.290 51.510 1413.610 51.570 ;
        RECT 1431.230 51.510 1431.550 51.570 ;
        RECT 1449.170 51.510 1449.490 51.570 ;
        RECT 1466.650 51.510 1466.970 51.570 ;
        RECT 1484.590 51.510 1484.910 51.570 ;
        RECT 1502.530 51.510 1502.850 51.570 ;
        RECT 1520.470 51.510 1520.790 51.570 ;
        RECT 1538.410 51.510 1538.730 51.570 ;
        RECT 1555.890 51.510 1556.210 51.570 ;
        RECT 1573.830 51.510 1574.150 51.570 ;
        RECT 1591.770 51.510 1592.090 51.570 ;
        RECT 1609.710 51.510 1610.030 51.570 ;
        RECT 1627.650 51.510 1627.970 51.570 ;
        RECT 1645.130 51.510 1645.450 51.570 ;
        RECT 1663.070 51.510 1663.390 51.570 ;
        RECT 1681.010 51.510 1681.330 51.570 ;
        RECT 1698.950 51.510 1699.270 51.570 ;
        RECT 1716.430 51.510 1716.750 51.570 ;
        RECT 1734.370 51.510 1734.690 51.570 ;
        RECT 1752.310 51.510 1752.630 51.570 ;
        RECT 1770.250 51.510 1770.570 51.570 ;
        RECT 1788.190 51.510 1788.510 51.570 ;
        RECT 1805.670 51.510 1805.990 51.570 ;
        RECT 1823.610 51.510 1823.930 51.570 ;
        RECT 1841.550 51.510 1841.870 51.570 ;
        RECT 1859.490 51.510 1859.810 51.570 ;
        RECT 1877.430 51.510 1877.750 51.570 ;
        RECT 1894.910 51.510 1895.230 51.570 ;
        RECT 1912.850 51.510 1913.170 51.570 ;
        RECT 1930.790 51.510 1931.110 51.570 ;
        RECT 1948.730 51.510 1949.050 51.570 ;
        RECT 1966.210 51.510 1966.530 51.570 ;
        RECT 1984.150 51.510 1984.470 51.570 ;
        RECT 2002.090 51.510 2002.410 51.570 ;
        RECT 2020.030 51.510 2020.350 51.570 ;
        RECT 2037.970 51.510 2038.290 51.570 ;
        RECT 2055.450 51.510 2055.770 51.570 ;
        RECT 2073.390 51.510 2073.710 51.570 ;
        RECT 2091.330 51.510 2091.650 51.570 ;
        RECT 2109.270 51.510 2109.590 51.570 ;
        RECT 2127.210 51.510 2127.530 51.570 ;
        RECT 2144.690 51.510 2145.010 51.570 ;
        RECT 2162.630 51.510 2162.950 51.570 ;
        RECT 2180.570 51.510 2180.890 51.570 ;
        RECT 2198.510 51.510 2198.830 51.570 ;
        RECT 2215.990 51.510 2216.310 51.570 ;
        RECT 2233.930 51.510 2234.250 51.570 ;
        RECT 2251.870 51.510 2252.190 51.570 ;
        RECT 2269.810 51.510 2270.130 51.570 ;
        RECT 2287.750 51.510 2288.070 51.570 ;
        RECT 2305.230 51.510 2305.550 51.570 ;
        RECT 2323.170 51.510 2323.490 51.570 ;
        RECT 2341.110 51.510 2341.430 51.570 ;
        RECT 2359.050 51.510 2359.370 51.570 ;
        RECT 2376.990 51.510 2377.310 51.570 ;
        RECT 2394.470 51.510 2394.790 51.570 ;
        RECT 2412.410 51.510 2412.730 51.570 ;
        RECT 2430.350 51.510 2430.670 51.570 ;
        RECT 2448.290 51.510 2448.610 51.570 ;
        RECT 2465.770 51.510 2466.090 51.570 ;
        RECT 2483.710 51.510 2484.030 51.570 ;
        RECT 2501.650 51.510 2501.970 51.570 ;
        RECT 2519.590 51.510 2519.910 51.570 ;
        RECT 2537.530 51.510 2537.850 51.570 ;
        RECT 2555.010 51.510 2555.330 51.570 ;
        RECT 2572.950 51.510 2573.270 51.570 ;
        RECT 2590.890 51.510 2591.210 51.570 ;
        RECT 2608.830 51.510 2609.150 51.570 ;
        RECT 2626.770 51.510 2627.090 51.570 ;
        RECT 2644.250 51.510 2644.570 51.570 ;
        RECT 2662.190 51.510 2662.510 51.570 ;
        RECT 2680.130 51.510 2680.450 51.570 ;
        RECT 2698.070 51.510 2698.390 51.570 ;
        RECT 2715.550 51.510 2715.870 51.570 ;
        RECT 2733.490 51.510 2733.810 51.570 ;
        RECT 2751.430 51.510 2751.750 51.570 ;
        RECT 2769.370 51.510 2769.690 51.570 ;
        RECT 2787.310 51.510 2787.630 51.570 ;
        RECT 2804.790 51.510 2805.110 51.570 ;
        RECT 2822.730 51.510 2823.050 51.570 ;
        RECT 2840.670 51.510 2840.990 51.570 ;
        RECT 2858.610 51.510 2858.930 51.570 ;
        RECT 2876.550 51.510 2876.870 51.570 ;
        RECT 2894.030 51.510 2894.350 51.570 ;
        RECT 2911.970 51.510 2912.290 51.570 ;
        RECT 2929.910 51.510 2930.230 51.570 ;
        RECT 2947.850 51.510 2948.170 51.570 ;
      LAYER via ;
        RECT 681.920 51.510 682.180 51.770 ;
        RECT 696.640 51.510 696.900 51.770 ;
        RECT 699.860 51.510 700.120 51.770 ;
        RECT 717.340 51.510 717.600 51.770 ;
        RECT 735.280 51.510 735.540 51.770 ;
        RECT 753.220 51.510 753.480 51.770 ;
        RECT 771.160 51.510 771.420 51.770 ;
        RECT 789.100 51.510 789.360 51.770 ;
        RECT 806.580 51.510 806.840 51.770 ;
        RECT 824.520 51.510 824.780 51.770 ;
        RECT 842.460 51.510 842.720 51.770 ;
        RECT 860.400 51.510 860.660 51.770 ;
        RECT 878.340 51.510 878.600 51.770 ;
        RECT 895.820 51.510 896.080 51.770 ;
        RECT 913.760 51.510 914.020 51.770 ;
        RECT 931.700 51.510 931.960 51.770 ;
        RECT 949.640 51.510 949.900 51.770 ;
        RECT 967.120 51.510 967.380 51.770 ;
        RECT 985.060 51.510 985.320 51.770 ;
        RECT 1003.000 51.510 1003.260 51.770 ;
        RECT 1020.940 51.510 1021.200 51.770 ;
        RECT 1038.880 51.510 1039.140 51.770 ;
        RECT 1056.360 51.510 1056.620 51.770 ;
        RECT 1074.300 51.510 1074.560 51.770 ;
        RECT 1092.240 51.510 1092.500 51.770 ;
        RECT 1110.180 51.510 1110.440 51.770 ;
        RECT 1128.120 51.510 1128.380 51.770 ;
        RECT 1145.600 51.510 1145.860 51.770 ;
        RECT 1163.540 51.510 1163.800 51.770 ;
        RECT 1181.480 51.510 1181.740 51.770 ;
        RECT 1199.420 51.510 1199.680 51.770 ;
        RECT 1216.900 51.510 1217.160 51.770 ;
        RECT 1234.840 51.510 1235.100 51.770 ;
        RECT 1252.780 51.510 1253.040 51.770 ;
        RECT 1270.720 51.510 1270.980 51.770 ;
        RECT 1288.660 51.510 1288.920 51.770 ;
        RECT 1306.140 51.510 1306.400 51.770 ;
        RECT 1324.080 51.510 1324.340 51.770 ;
        RECT 1342.020 51.510 1342.280 51.770 ;
        RECT 1359.960 51.510 1360.220 51.770 ;
        RECT 1377.900 51.510 1378.160 51.770 ;
        RECT 1395.380 51.510 1395.640 51.770 ;
        RECT 1413.320 51.510 1413.580 51.770 ;
        RECT 1431.260 51.510 1431.520 51.770 ;
        RECT 1449.200 51.510 1449.460 51.770 ;
        RECT 1466.680 51.510 1466.940 51.770 ;
        RECT 1484.620 51.510 1484.880 51.770 ;
        RECT 1502.560 51.510 1502.820 51.770 ;
        RECT 1520.500 51.510 1520.760 51.770 ;
        RECT 1538.440 51.510 1538.700 51.770 ;
        RECT 1555.920 51.510 1556.180 51.770 ;
        RECT 1573.860 51.510 1574.120 51.770 ;
        RECT 1591.800 51.510 1592.060 51.770 ;
        RECT 1609.740 51.510 1610.000 51.770 ;
        RECT 1627.680 51.510 1627.940 51.770 ;
        RECT 1645.160 51.510 1645.420 51.770 ;
        RECT 1663.100 51.510 1663.360 51.770 ;
        RECT 1681.040 51.510 1681.300 51.770 ;
        RECT 1698.980 51.510 1699.240 51.770 ;
        RECT 1716.460 51.510 1716.720 51.770 ;
        RECT 1734.400 51.510 1734.660 51.770 ;
        RECT 1752.340 51.510 1752.600 51.770 ;
        RECT 1770.280 51.510 1770.540 51.770 ;
        RECT 1788.220 51.510 1788.480 51.770 ;
        RECT 1805.700 51.510 1805.960 51.770 ;
        RECT 1823.640 51.510 1823.900 51.770 ;
        RECT 1841.580 51.510 1841.840 51.770 ;
        RECT 1859.520 51.510 1859.780 51.770 ;
        RECT 1877.460 51.510 1877.720 51.770 ;
        RECT 1894.940 51.510 1895.200 51.770 ;
        RECT 1912.880 51.510 1913.140 51.770 ;
        RECT 1930.820 51.510 1931.080 51.770 ;
        RECT 1948.760 51.510 1949.020 51.770 ;
        RECT 1966.240 51.510 1966.500 51.770 ;
        RECT 1984.180 51.510 1984.440 51.770 ;
        RECT 2002.120 51.510 2002.380 51.770 ;
        RECT 2020.060 51.510 2020.320 51.770 ;
        RECT 2038.000 51.510 2038.260 51.770 ;
        RECT 2055.480 51.510 2055.740 51.770 ;
        RECT 2073.420 51.510 2073.680 51.770 ;
        RECT 2091.360 51.510 2091.620 51.770 ;
        RECT 2109.300 51.510 2109.560 51.770 ;
        RECT 2127.240 51.510 2127.500 51.770 ;
        RECT 2144.720 51.510 2144.980 51.770 ;
        RECT 2162.660 51.510 2162.920 51.770 ;
        RECT 2180.600 51.510 2180.860 51.770 ;
        RECT 2198.540 51.510 2198.800 51.770 ;
        RECT 2216.020 51.510 2216.280 51.770 ;
        RECT 2233.960 51.510 2234.220 51.770 ;
        RECT 2251.900 51.510 2252.160 51.770 ;
        RECT 2269.840 51.510 2270.100 51.770 ;
        RECT 2287.780 51.510 2288.040 51.770 ;
        RECT 2305.260 51.510 2305.520 51.770 ;
        RECT 2323.200 51.510 2323.460 51.770 ;
        RECT 2341.140 51.510 2341.400 51.770 ;
        RECT 2359.080 51.510 2359.340 51.770 ;
        RECT 2377.020 51.510 2377.280 51.770 ;
        RECT 2394.500 51.510 2394.760 51.770 ;
        RECT 2412.440 51.510 2412.700 51.770 ;
        RECT 2430.380 51.510 2430.640 51.770 ;
        RECT 2448.320 51.510 2448.580 51.770 ;
        RECT 2465.800 51.510 2466.060 51.770 ;
        RECT 2483.740 51.510 2484.000 51.770 ;
        RECT 2501.680 51.510 2501.940 51.770 ;
        RECT 2519.620 51.510 2519.880 51.770 ;
        RECT 2537.560 51.510 2537.820 51.770 ;
        RECT 2555.040 51.510 2555.300 51.770 ;
        RECT 2572.980 51.510 2573.240 51.770 ;
        RECT 2590.920 51.510 2591.180 51.770 ;
        RECT 2608.860 51.510 2609.120 51.770 ;
        RECT 2626.800 51.510 2627.060 51.770 ;
        RECT 2644.280 51.510 2644.540 51.770 ;
        RECT 2662.220 51.510 2662.480 51.770 ;
        RECT 2680.160 51.510 2680.420 51.770 ;
        RECT 2698.100 51.510 2698.360 51.770 ;
        RECT 2715.580 51.510 2715.840 51.770 ;
        RECT 2733.520 51.510 2733.780 51.770 ;
        RECT 2751.460 51.510 2751.720 51.770 ;
        RECT 2769.400 51.510 2769.660 51.770 ;
        RECT 2787.340 51.510 2787.600 51.770 ;
        RECT 2804.820 51.510 2805.080 51.770 ;
        RECT 2822.760 51.510 2823.020 51.770 ;
        RECT 2840.700 51.510 2840.960 51.770 ;
        RECT 2858.640 51.510 2858.900 51.770 ;
        RECT 2876.580 51.510 2876.840 51.770 ;
        RECT 2894.060 51.510 2894.320 51.770 ;
        RECT 2912.000 51.510 2912.260 51.770 ;
        RECT 2929.940 51.510 2930.200 51.770 ;
        RECT 2947.880 51.510 2948.140 51.770 ;
      LAYER met2 ;
        RECT 696.700 51.800 696.840 54.000 ;
        RECT 681.920 51.480 682.180 51.800 ;
        RECT 696.640 51.480 696.900 51.800 ;
        RECT 699.860 51.480 700.120 51.800 ;
        RECT 717.340 51.480 717.600 51.800 ;
        RECT 735.280 51.480 735.540 51.800 ;
        RECT 753.220 51.480 753.480 51.800 ;
        RECT 771.160 51.480 771.420 51.800 ;
        RECT 789.100 51.480 789.360 51.800 ;
        RECT 806.580 51.480 806.840 51.800 ;
        RECT 824.520 51.480 824.780 51.800 ;
        RECT 842.460 51.480 842.720 51.800 ;
        RECT 860.400 51.480 860.660 51.800 ;
        RECT 878.340 51.480 878.600 51.800 ;
        RECT 895.820 51.480 896.080 51.800 ;
        RECT 913.760 51.480 914.020 51.800 ;
        RECT 931.700 51.480 931.960 51.800 ;
        RECT 949.640 51.480 949.900 51.800 ;
        RECT 967.120 51.480 967.380 51.800 ;
        RECT 985.060 51.480 985.320 51.800 ;
        RECT 1003.000 51.480 1003.260 51.800 ;
        RECT 1020.940 51.480 1021.200 51.800 ;
        RECT 1038.880 51.480 1039.140 51.800 ;
        RECT 1056.360 51.480 1056.620 51.800 ;
        RECT 1074.300 51.480 1074.560 51.800 ;
        RECT 1092.240 51.480 1092.500 51.800 ;
        RECT 1110.180 51.480 1110.440 51.800 ;
        RECT 1128.120 51.480 1128.380 51.800 ;
        RECT 1145.600 51.480 1145.860 51.800 ;
        RECT 1163.540 51.480 1163.800 51.800 ;
        RECT 1181.480 51.480 1181.740 51.800 ;
        RECT 1199.420 51.480 1199.680 51.800 ;
        RECT 1216.900 51.480 1217.160 51.800 ;
        RECT 1234.840 51.480 1235.100 51.800 ;
        RECT 1252.780 51.480 1253.040 51.800 ;
        RECT 1270.720 51.480 1270.980 51.800 ;
        RECT 1288.660 51.480 1288.920 51.800 ;
        RECT 1306.140 51.480 1306.400 51.800 ;
        RECT 1324.080 51.480 1324.340 51.800 ;
        RECT 1342.020 51.480 1342.280 51.800 ;
        RECT 1359.960 51.480 1360.220 51.800 ;
        RECT 1377.900 51.480 1378.160 51.800 ;
        RECT 1395.380 51.480 1395.640 51.800 ;
        RECT 1413.320 51.480 1413.580 51.800 ;
        RECT 1431.260 51.480 1431.520 51.800 ;
        RECT 1449.200 51.480 1449.460 51.800 ;
        RECT 1466.680 51.480 1466.940 51.800 ;
        RECT 1484.620 51.480 1484.880 51.800 ;
        RECT 1502.560 51.480 1502.820 51.800 ;
        RECT 1520.500 51.480 1520.760 51.800 ;
        RECT 1538.440 51.480 1538.700 51.800 ;
        RECT 1555.920 51.480 1556.180 51.800 ;
        RECT 1573.860 51.480 1574.120 51.800 ;
        RECT 1591.800 51.480 1592.060 51.800 ;
        RECT 1609.740 51.480 1610.000 51.800 ;
        RECT 1627.680 51.480 1627.940 51.800 ;
        RECT 1645.160 51.480 1645.420 51.800 ;
        RECT 1663.100 51.480 1663.360 51.800 ;
        RECT 1681.040 51.480 1681.300 51.800 ;
        RECT 1698.980 51.480 1699.240 51.800 ;
        RECT 1716.460 51.480 1716.720 51.800 ;
        RECT 1734.400 51.480 1734.660 51.800 ;
        RECT 1752.340 51.480 1752.600 51.800 ;
        RECT 1770.280 51.480 1770.540 51.800 ;
        RECT 1788.220 51.480 1788.480 51.800 ;
        RECT 1805.700 51.480 1805.960 51.800 ;
        RECT 1823.640 51.480 1823.900 51.800 ;
        RECT 1841.580 51.480 1841.840 51.800 ;
        RECT 1859.520 51.480 1859.780 51.800 ;
        RECT 1877.460 51.480 1877.720 51.800 ;
        RECT 1894.940 51.480 1895.200 51.800 ;
        RECT 1912.880 51.480 1913.140 51.800 ;
        RECT 1930.820 51.480 1931.080 51.800 ;
        RECT 1948.760 51.480 1949.020 51.800 ;
        RECT 1966.240 51.480 1966.500 51.800 ;
        RECT 1984.180 51.480 1984.440 51.800 ;
        RECT 2002.120 51.480 2002.380 51.800 ;
        RECT 2020.060 51.480 2020.320 51.800 ;
        RECT 2038.000 51.480 2038.260 51.800 ;
        RECT 2055.480 51.480 2055.740 51.800 ;
        RECT 2073.420 51.480 2073.680 51.800 ;
        RECT 2091.360 51.480 2091.620 51.800 ;
        RECT 2109.300 51.480 2109.560 51.800 ;
        RECT 2127.240 51.480 2127.500 51.800 ;
        RECT 2144.720 51.480 2144.980 51.800 ;
        RECT 2162.660 51.480 2162.920 51.800 ;
        RECT 2180.600 51.480 2180.860 51.800 ;
        RECT 2198.540 51.480 2198.800 51.800 ;
        RECT 2216.020 51.480 2216.280 51.800 ;
        RECT 2233.960 51.480 2234.220 51.800 ;
        RECT 2251.900 51.480 2252.160 51.800 ;
        RECT 2269.840 51.480 2270.100 51.800 ;
        RECT 2287.780 51.480 2288.040 51.800 ;
        RECT 2305.260 51.480 2305.520 51.800 ;
        RECT 2323.200 51.480 2323.460 51.800 ;
        RECT 2341.140 51.480 2341.400 51.800 ;
        RECT 2359.080 51.480 2359.340 51.800 ;
        RECT 2377.020 51.480 2377.280 51.800 ;
        RECT 2394.500 51.480 2394.760 51.800 ;
        RECT 2412.440 51.480 2412.700 51.800 ;
        RECT 2430.380 51.480 2430.640 51.800 ;
        RECT 2448.320 51.480 2448.580 51.800 ;
        RECT 2465.800 51.480 2466.060 51.800 ;
        RECT 2483.740 51.480 2484.000 51.800 ;
        RECT 2501.680 51.480 2501.940 51.800 ;
        RECT 2519.620 51.480 2519.880 51.800 ;
        RECT 2537.560 51.480 2537.820 51.800 ;
        RECT 2555.040 51.480 2555.300 51.800 ;
        RECT 2572.980 51.480 2573.240 51.800 ;
        RECT 2590.920 51.480 2591.180 51.800 ;
        RECT 2608.860 51.480 2609.120 51.800 ;
        RECT 2626.800 51.480 2627.060 51.800 ;
        RECT 2644.280 51.480 2644.540 51.800 ;
        RECT 2662.220 51.480 2662.480 51.800 ;
        RECT 2680.160 51.480 2680.420 51.800 ;
        RECT 2698.100 51.480 2698.360 51.800 ;
        RECT 2715.580 51.480 2715.840 51.800 ;
        RECT 2733.520 51.480 2733.780 51.800 ;
        RECT 2751.460 51.480 2751.720 51.800 ;
        RECT 2769.400 51.480 2769.660 51.800 ;
        RECT 2787.340 51.480 2787.600 51.800 ;
        RECT 2804.820 51.480 2805.080 51.800 ;
        RECT 2822.760 51.480 2823.020 51.800 ;
        RECT 2840.700 51.480 2840.960 51.800 ;
        RECT 2858.640 51.480 2858.900 51.800 ;
        RECT 2876.580 51.480 2876.840 51.800 ;
        RECT 2894.060 51.480 2894.320 51.800 ;
        RECT 2912.000 51.480 2912.260 51.800 ;
        RECT 2929.940 51.480 2930.200 51.800 ;
        RECT 2947.880 51.480 2948.140 51.800 ;
        RECT 681.980 41.530 682.120 51.480 ;
        RECT 699.920 41.530 700.060 51.480 ;
        RECT 717.400 41.530 717.540 51.480 ;
        RECT 735.340 41.530 735.480 51.480 ;
        RECT 753.280 41.530 753.420 51.480 ;
        RECT 771.220 41.530 771.360 51.480 ;
        RECT 789.160 41.530 789.300 51.480 ;
        RECT 806.640 41.530 806.780 51.480 ;
        RECT 824.580 41.530 824.720 51.480 ;
        RECT 842.520 41.530 842.660 51.480 ;
        RECT 860.460 41.530 860.600 51.480 ;
        RECT 878.400 41.530 878.540 51.480 ;
        RECT 895.880 41.530 896.020 51.480 ;
        RECT 913.820 41.530 913.960 51.480 ;
        RECT 931.760 41.530 931.900 51.480 ;
        RECT 949.700 41.530 949.840 51.480 ;
        RECT 967.180 41.530 967.320 51.480 ;
        RECT 985.120 41.530 985.260 51.480 ;
        RECT 1003.060 41.530 1003.200 51.480 ;
        RECT 1021.000 41.530 1021.140 51.480 ;
        RECT 1038.940 41.530 1039.080 51.480 ;
        RECT 1056.420 41.530 1056.560 51.480 ;
        RECT 1074.360 41.530 1074.500 51.480 ;
        RECT 1092.300 41.530 1092.440 51.480 ;
        RECT 1110.240 41.530 1110.380 51.480 ;
        RECT 1128.180 41.530 1128.320 51.480 ;
        RECT 1145.660 41.530 1145.800 51.480 ;
        RECT 1163.600 41.530 1163.740 51.480 ;
        RECT 1181.540 41.530 1181.680 51.480 ;
        RECT 1199.480 41.530 1199.620 51.480 ;
        RECT 1216.960 41.530 1217.100 51.480 ;
        RECT 1234.900 41.530 1235.040 51.480 ;
        RECT 1252.840 41.530 1252.980 51.480 ;
        RECT 1270.780 41.530 1270.920 51.480 ;
        RECT 1288.720 41.530 1288.860 51.480 ;
        RECT 1306.200 41.530 1306.340 51.480 ;
        RECT 1324.140 41.530 1324.280 51.480 ;
        RECT 1342.080 41.530 1342.220 51.480 ;
        RECT 1360.020 41.530 1360.160 51.480 ;
        RECT 1377.960 41.530 1378.100 51.480 ;
        RECT 1395.440 41.530 1395.580 51.480 ;
        RECT 1413.380 41.530 1413.520 51.480 ;
        RECT 1431.320 41.530 1431.460 51.480 ;
        RECT 1449.260 41.530 1449.400 51.480 ;
        RECT 1466.740 41.530 1466.880 51.480 ;
        RECT 1484.680 41.530 1484.820 51.480 ;
        RECT 1502.620 41.530 1502.760 51.480 ;
        RECT 1520.560 41.530 1520.700 51.480 ;
        RECT 1538.500 41.530 1538.640 51.480 ;
        RECT 1555.980 41.530 1556.120 51.480 ;
        RECT 1573.920 41.530 1574.060 51.480 ;
        RECT 1591.860 41.530 1592.000 51.480 ;
        RECT 1609.800 41.530 1609.940 51.480 ;
        RECT 1627.740 41.530 1627.880 51.480 ;
        RECT 1645.220 41.530 1645.360 51.480 ;
        RECT 1663.160 41.530 1663.300 51.480 ;
        RECT 1681.100 41.530 1681.240 51.480 ;
        RECT 1699.040 41.530 1699.180 51.480 ;
        RECT 1716.520 41.530 1716.660 51.480 ;
        RECT 1734.460 41.530 1734.600 51.480 ;
        RECT 1752.400 41.530 1752.540 51.480 ;
        RECT 1770.340 41.530 1770.480 51.480 ;
        RECT 1788.280 41.530 1788.420 51.480 ;
        RECT 1805.760 41.530 1805.900 51.480 ;
        RECT 1823.700 41.530 1823.840 51.480 ;
        RECT 1841.640 41.530 1841.780 51.480 ;
        RECT 1859.580 41.530 1859.720 51.480 ;
        RECT 1877.520 41.530 1877.660 51.480 ;
        RECT 1895.000 41.530 1895.140 51.480 ;
        RECT 1912.940 41.530 1913.080 51.480 ;
        RECT 1930.880 41.530 1931.020 51.480 ;
        RECT 1948.820 41.530 1948.960 51.480 ;
        RECT 1966.300 41.530 1966.440 51.480 ;
        RECT 1984.240 41.530 1984.380 51.480 ;
        RECT 2002.180 41.530 2002.320 51.480 ;
        RECT 2020.120 41.530 2020.260 51.480 ;
        RECT 2038.060 41.530 2038.200 51.480 ;
        RECT 2055.540 41.530 2055.680 51.480 ;
        RECT 2073.480 41.530 2073.620 51.480 ;
        RECT 2091.420 41.530 2091.560 51.480 ;
        RECT 2109.360 41.530 2109.500 51.480 ;
        RECT 2127.300 41.530 2127.440 51.480 ;
        RECT 2144.780 41.530 2144.920 51.480 ;
        RECT 2162.720 41.530 2162.860 51.480 ;
        RECT 2180.660 41.530 2180.800 51.480 ;
        RECT 2198.600 41.530 2198.740 51.480 ;
        RECT 2216.080 41.530 2216.220 51.480 ;
        RECT 2234.020 41.530 2234.160 51.480 ;
        RECT 2251.960 41.530 2252.100 51.480 ;
        RECT 2269.900 41.530 2270.040 51.480 ;
        RECT 2287.840 41.530 2287.980 51.480 ;
        RECT 2305.320 41.530 2305.460 51.480 ;
        RECT 2323.260 41.530 2323.400 51.480 ;
        RECT 2341.200 41.530 2341.340 51.480 ;
        RECT 2359.140 41.530 2359.280 51.480 ;
        RECT 2377.080 41.530 2377.220 51.480 ;
        RECT 2394.560 41.530 2394.700 51.480 ;
        RECT 2412.500 41.530 2412.640 51.480 ;
        RECT 2430.440 41.530 2430.580 51.480 ;
        RECT 2448.380 41.530 2448.520 51.480 ;
        RECT 2465.860 41.530 2466.000 51.480 ;
        RECT 2483.800 41.530 2483.940 51.480 ;
        RECT 2501.740 41.530 2501.880 51.480 ;
        RECT 2519.680 41.530 2519.820 51.480 ;
        RECT 2537.620 41.530 2537.760 51.480 ;
        RECT 2555.100 41.530 2555.240 51.480 ;
        RECT 2573.040 41.530 2573.180 51.480 ;
        RECT 2590.980 41.530 2591.120 51.480 ;
        RECT 2608.920 41.530 2609.060 51.480 ;
        RECT 2626.860 41.530 2627.000 51.480 ;
        RECT 2644.340 41.530 2644.480 51.480 ;
        RECT 2662.280 41.530 2662.420 51.480 ;
        RECT 2680.220 41.530 2680.360 51.480 ;
        RECT 2698.160 41.530 2698.300 51.480 ;
        RECT 2715.640 41.530 2715.780 51.480 ;
        RECT 2733.580 41.530 2733.720 51.480 ;
        RECT 2751.520 41.530 2751.660 51.480 ;
        RECT 2769.460 41.530 2769.600 51.480 ;
        RECT 2787.400 41.530 2787.540 51.480 ;
        RECT 2804.880 41.530 2805.020 51.480 ;
        RECT 2822.820 41.530 2822.960 51.480 ;
        RECT 2840.760 41.530 2840.900 51.480 ;
        RECT 2858.700 41.530 2858.840 51.480 ;
        RECT 2876.640 41.530 2876.780 51.480 ;
        RECT 2894.120 41.530 2894.260 51.480 ;
        RECT 2912.060 41.530 2912.200 51.480 ;
        RECT 2930.000 41.530 2930.140 51.480 ;
        RECT 2947.940 41.530 2948.080 51.480 ;
        RECT 681.910 37.530 682.190 41.530 ;
        RECT 699.850 37.530 700.130 41.530 ;
        RECT 717.330 37.530 717.610 41.530 ;
        RECT 735.270 37.530 735.550 41.530 ;
        RECT 753.210 37.530 753.490 41.530 ;
        RECT 771.150 37.530 771.430 41.530 ;
        RECT 789.090 37.530 789.370 41.530 ;
        RECT 806.570 37.530 806.850 41.530 ;
        RECT 824.510 37.530 824.790 41.530 ;
        RECT 842.450 37.530 842.730 41.530 ;
        RECT 860.390 37.530 860.670 41.530 ;
        RECT 878.330 37.530 878.610 41.530 ;
        RECT 895.810 37.530 896.090 41.530 ;
        RECT 913.750 37.530 914.030 41.530 ;
        RECT 931.690 37.530 931.970 41.530 ;
        RECT 949.630 37.530 949.910 41.530 ;
        RECT 967.110 37.530 967.390 41.530 ;
        RECT 985.050 37.530 985.330 41.530 ;
        RECT 1002.990 37.530 1003.270 41.530 ;
        RECT 1020.930 37.530 1021.210 41.530 ;
        RECT 1038.870 37.530 1039.150 41.530 ;
        RECT 1056.350 37.530 1056.630 41.530 ;
        RECT 1074.290 37.530 1074.570 41.530 ;
        RECT 1092.230 37.530 1092.510 41.530 ;
        RECT 1110.170 37.530 1110.450 41.530 ;
        RECT 1128.110 37.530 1128.390 41.530 ;
        RECT 1145.590 37.530 1145.870 41.530 ;
        RECT 1163.530 37.530 1163.810 41.530 ;
        RECT 1181.470 37.530 1181.750 41.530 ;
        RECT 1199.410 37.530 1199.690 41.530 ;
        RECT 1216.890 37.530 1217.170 41.530 ;
        RECT 1234.830 37.530 1235.110 41.530 ;
        RECT 1252.770 37.530 1253.050 41.530 ;
        RECT 1270.710 37.530 1270.990 41.530 ;
        RECT 1288.650 37.530 1288.930 41.530 ;
        RECT 1306.130 37.530 1306.410 41.530 ;
        RECT 1324.070 37.530 1324.350 41.530 ;
        RECT 1342.010 37.530 1342.290 41.530 ;
        RECT 1359.950 37.530 1360.230 41.530 ;
        RECT 1377.890 37.530 1378.170 41.530 ;
        RECT 1395.370 37.530 1395.650 41.530 ;
        RECT 1413.310 37.530 1413.590 41.530 ;
        RECT 1431.250 37.530 1431.530 41.530 ;
        RECT 1449.190 37.530 1449.470 41.530 ;
        RECT 1466.670 37.530 1466.950 41.530 ;
        RECT 1484.610 37.530 1484.890 41.530 ;
        RECT 1502.550 37.530 1502.830 41.530 ;
        RECT 1520.490 37.530 1520.770 41.530 ;
        RECT 1538.430 37.530 1538.710 41.530 ;
        RECT 1555.910 37.530 1556.190 41.530 ;
        RECT 1573.850 37.530 1574.130 41.530 ;
        RECT 1591.790 37.530 1592.070 41.530 ;
        RECT 1609.730 37.530 1610.010 41.530 ;
        RECT 1627.670 37.530 1627.950 41.530 ;
        RECT 1645.150 37.530 1645.430 41.530 ;
        RECT 1663.090 37.530 1663.370 41.530 ;
        RECT 1681.030 37.530 1681.310 41.530 ;
        RECT 1698.970 37.530 1699.250 41.530 ;
        RECT 1716.450 37.530 1716.730 41.530 ;
        RECT 1734.390 37.530 1734.670 41.530 ;
        RECT 1752.330 37.530 1752.610 41.530 ;
        RECT 1770.270 37.530 1770.550 41.530 ;
        RECT 1788.210 37.530 1788.490 41.530 ;
        RECT 1805.690 37.530 1805.970 41.530 ;
        RECT 1823.630 37.530 1823.910 41.530 ;
        RECT 1841.570 37.530 1841.850 41.530 ;
        RECT 1859.510 37.530 1859.790 41.530 ;
        RECT 1877.450 37.530 1877.730 41.530 ;
        RECT 1894.930 37.530 1895.210 41.530 ;
        RECT 1912.870 37.530 1913.150 41.530 ;
        RECT 1930.810 37.530 1931.090 41.530 ;
        RECT 1948.750 37.530 1949.030 41.530 ;
        RECT 1966.230 37.530 1966.510 41.530 ;
        RECT 1984.170 37.530 1984.450 41.530 ;
        RECT 2002.110 37.530 2002.390 41.530 ;
        RECT 2020.050 37.530 2020.330 41.530 ;
        RECT 2037.990 37.530 2038.270 41.530 ;
        RECT 2055.470 37.530 2055.750 41.530 ;
        RECT 2073.410 37.530 2073.690 41.530 ;
        RECT 2091.350 37.530 2091.630 41.530 ;
        RECT 2109.290 37.530 2109.570 41.530 ;
        RECT 2127.230 37.530 2127.510 41.530 ;
        RECT 2144.710 37.530 2144.990 41.530 ;
        RECT 2162.650 37.530 2162.930 41.530 ;
        RECT 2180.590 37.530 2180.870 41.530 ;
        RECT 2198.530 37.530 2198.810 41.530 ;
        RECT 2216.010 37.530 2216.290 41.530 ;
        RECT 2233.950 37.530 2234.230 41.530 ;
        RECT 2251.890 37.530 2252.170 41.530 ;
        RECT 2269.830 37.530 2270.110 41.530 ;
        RECT 2287.770 37.530 2288.050 41.530 ;
        RECT 2305.250 37.530 2305.530 41.530 ;
        RECT 2323.190 37.530 2323.470 41.530 ;
        RECT 2341.130 37.530 2341.410 41.530 ;
        RECT 2359.070 37.530 2359.350 41.530 ;
        RECT 2377.010 37.530 2377.290 41.530 ;
        RECT 2394.490 37.530 2394.770 41.530 ;
        RECT 2412.430 37.530 2412.710 41.530 ;
        RECT 2430.370 37.530 2430.650 41.530 ;
        RECT 2448.310 37.530 2448.590 41.530 ;
        RECT 2465.790 37.530 2466.070 41.530 ;
        RECT 2483.730 37.530 2484.010 41.530 ;
        RECT 2501.670 37.530 2501.950 41.530 ;
        RECT 2519.610 37.530 2519.890 41.530 ;
        RECT 2537.550 37.530 2537.830 41.530 ;
        RECT 2555.030 37.530 2555.310 41.530 ;
        RECT 2572.970 37.530 2573.250 41.530 ;
        RECT 2590.910 37.530 2591.190 41.530 ;
        RECT 2608.850 37.530 2609.130 41.530 ;
        RECT 2626.790 37.530 2627.070 41.530 ;
        RECT 2644.270 37.530 2644.550 41.530 ;
        RECT 2662.210 37.530 2662.490 41.530 ;
        RECT 2680.150 37.530 2680.430 41.530 ;
        RECT 2698.090 37.530 2698.370 41.530 ;
        RECT 2715.570 37.530 2715.850 41.530 ;
        RECT 2733.510 37.530 2733.790 41.530 ;
        RECT 2751.450 37.530 2751.730 41.530 ;
        RECT 2769.390 37.530 2769.670 41.530 ;
        RECT 2787.330 37.530 2787.610 41.530 ;
        RECT 2804.810 37.530 2805.090 41.530 ;
        RECT 2822.750 37.530 2823.030 41.530 ;
        RECT 2840.690 37.530 2840.970 41.530 ;
        RECT 2858.630 37.530 2858.910 41.530 ;
        RECT 2876.570 37.530 2876.850 41.530 ;
        RECT 2894.050 37.530 2894.330 41.530 ;
        RECT 2911.990 37.530 2912.270 41.530 ;
        RECT 2929.930 37.530 2930.210 41.530 ;
        RECT 2947.870 37.530 2948.150 41.530 ;
    END
  END la_data_out[0]
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 32.900 32.910 35.900 3561.830 ;
        RECT 46.900 28.210 49.900 3566.530 ;
        RECT 226.900 3540.740 229.900 3566.530 ;
        RECT 406.900 3540.740 409.900 3566.530 ;
        RECT 586.900 3540.740 589.900 3566.530 ;
        RECT 766.900 3540.740 769.900 3566.530 ;
        RECT 946.900 3540.740 949.900 3566.530 ;
        RECT 1126.900 3540.740 1129.900 3566.530 ;
        RECT 1306.900 3540.740 1309.900 3566.530 ;
        RECT 1486.900 3540.740 1489.900 3566.530 ;
        RECT 1666.900 3540.740 1669.900 3566.530 ;
        RECT 1846.900 3540.740 1849.900 3566.530 ;
        RECT 2026.900 3540.740 2029.900 3566.530 ;
        RECT 2206.900 3540.740 2209.900 3566.530 ;
        RECT 2386.900 3540.740 2389.900 3566.530 ;
        RECT 2566.900 3540.740 2569.900 3566.530 ;
        RECT 2746.900 3540.740 2749.900 3566.530 ;
        RECT 2926.900 3540.740 2929.900 3566.530 ;
        RECT 226.900 28.210 229.900 54.000 ;
        RECT 406.900 28.210 409.900 54.000 ;
        RECT 586.900 28.210 589.900 54.000 ;
        RECT 766.900 28.210 769.900 54.000 ;
        RECT 946.900 28.210 949.900 54.000 ;
        RECT 1126.900 28.210 1129.900 54.000 ;
        RECT 1306.900 28.210 1309.900 54.000 ;
        RECT 1486.900 28.210 1489.900 54.000 ;
        RECT 1666.900 28.210 1669.900 54.000 ;
        RECT 1846.900 28.210 1849.900 54.000 ;
        RECT 2026.900 28.210 2029.900 54.000 ;
        RECT 2206.900 28.210 2209.900 54.000 ;
        RECT 2386.900 28.210 2389.900 54.000 ;
        RECT 2566.900 28.210 2569.900 54.000 ;
        RECT 2746.900 28.210 2749.900 54.000 ;
        RECT 2926.900 28.210 2929.900 54.000 ;
        RECT 2969.480 32.910 2972.480 3561.830 ;
      LAYER M4M5_PR_C ;
        RECT 33.810 3560.540 34.990 3561.720 ;
        RECT 33.810 3558.940 34.990 3560.120 ;
        RECT 33.810 3468.620 34.990 3469.800 ;
        RECT 33.810 3467.020 34.990 3468.200 ;
        RECT 33.810 3288.620 34.990 3289.800 ;
        RECT 33.810 3287.020 34.990 3288.200 ;
        RECT 33.810 3108.620 34.990 3109.800 ;
        RECT 33.810 3107.020 34.990 3108.200 ;
        RECT 33.810 2928.620 34.990 2929.800 ;
        RECT 33.810 2927.020 34.990 2928.200 ;
        RECT 33.810 2748.620 34.990 2749.800 ;
        RECT 33.810 2747.020 34.990 2748.200 ;
        RECT 33.810 2568.620 34.990 2569.800 ;
        RECT 33.810 2567.020 34.990 2568.200 ;
        RECT 33.810 2388.620 34.990 2389.800 ;
        RECT 33.810 2387.020 34.990 2388.200 ;
        RECT 33.810 2208.620 34.990 2209.800 ;
        RECT 33.810 2207.020 34.990 2208.200 ;
        RECT 33.810 2028.620 34.990 2029.800 ;
        RECT 33.810 2027.020 34.990 2028.200 ;
        RECT 33.810 1848.620 34.990 1849.800 ;
        RECT 33.810 1847.020 34.990 1848.200 ;
        RECT 33.810 1668.620 34.990 1669.800 ;
        RECT 33.810 1667.020 34.990 1668.200 ;
        RECT 33.810 1488.620 34.990 1489.800 ;
        RECT 33.810 1487.020 34.990 1488.200 ;
        RECT 33.810 1308.620 34.990 1309.800 ;
        RECT 33.810 1307.020 34.990 1308.200 ;
        RECT 33.810 1128.620 34.990 1129.800 ;
        RECT 33.810 1127.020 34.990 1128.200 ;
        RECT 33.810 948.620 34.990 949.800 ;
        RECT 33.810 947.020 34.990 948.200 ;
        RECT 33.810 768.620 34.990 769.800 ;
        RECT 33.810 767.020 34.990 768.200 ;
        RECT 33.810 588.620 34.990 589.800 ;
        RECT 33.810 587.020 34.990 588.200 ;
        RECT 33.810 408.620 34.990 409.800 ;
        RECT 33.810 407.020 34.990 408.200 ;
        RECT 33.810 228.620 34.990 229.800 ;
        RECT 33.810 227.020 34.990 228.200 ;
        RECT 33.810 48.620 34.990 49.800 ;
        RECT 33.810 47.020 34.990 48.200 ;
        RECT 33.810 34.620 34.990 35.800 ;
        RECT 33.810 33.020 34.990 34.200 ;
        RECT 47.810 3560.540 48.990 3561.720 ;
        RECT 47.810 3558.940 48.990 3560.120 ;
        RECT 227.810 3560.540 228.990 3561.720 ;
        RECT 227.810 3558.940 228.990 3560.120 ;
        RECT 407.810 3560.540 408.990 3561.720 ;
        RECT 407.810 3558.940 408.990 3560.120 ;
        RECT 587.810 3560.540 588.990 3561.720 ;
        RECT 587.810 3558.940 588.990 3560.120 ;
        RECT 767.810 3560.540 768.990 3561.720 ;
        RECT 767.810 3558.940 768.990 3560.120 ;
        RECT 947.810 3560.540 948.990 3561.720 ;
        RECT 947.810 3558.940 948.990 3560.120 ;
        RECT 1127.810 3560.540 1128.990 3561.720 ;
        RECT 1127.810 3558.940 1128.990 3560.120 ;
        RECT 1307.810 3560.540 1308.990 3561.720 ;
        RECT 1307.810 3558.940 1308.990 3560.120 ;
        RECT 1487.810 3560.540 1488.990 3561.720 ;
        RECT 1487.810 3558.940 1488.990 3560.120 ;
        RECT 1667.810 3560.540 1668.990 3561.720 ;
        RECT 1667.810 3558.940 1668.990 3560.120 ;
        RECT 1847.810 3560.540 1848.990 3561.720 ;
        RECT 1847.810 3558.940 1848.990 3560.120 ;
        RECT 2027.810 3560.540 2028.990 3561.720 ;
        RECT 2027.810 3558.940 2028.990 3560.120 ;
        RECT 2207.810 3560.540 2208.990 3561.720 ;
        RECT 2207.810 3558.940 2208.990 3560.120 ;
        RECT 2387.810 3560.540 2388.990 3561.720 ;
        RECT 2387.810 3558.940 2388.990 3560.120 ;
        RECT 2567.810 3560.540 2568.990 3561.720 ;
        RECT 2567.810 3558.940 2568.990 3560.120 ;
        RECT 2747.810 3560.540 2748.990 3561.720 ;
        RECT 2747.810 3558.940 2748.990 3560.120 ;
        RECT 2927.810 3560.540 2928.990 3561.720 ;
        RECT 2927.810 3558.940 2928.990 3560.120 ;
        RECT 2970.390 3560.540 2971.570 3561.720 ;
        RECT 2970.390 3558.940 2971.570 3560.120 ;
        RECT 47.810 3468.620 48.990 3469.800 ;
        RECT 47.810 3467.020 48.990 3468.200 ;
        RECT 47.810 3288.620 48.990 3289.800 ;
        RECT 47.810 3287.020 48.990 3288.200 ;
        RECT 47.810 3108.620 48.990 3109.800 ;
        RECT 47.810 3107.020 48.990 3108.200 ;
        RECT 47.810 2928.620 48.990 2929.800 ;
        RECT 47.810 2927.020 48.990 2928.200 ;
        RECT 47.810 2748.620 48.990 2749.800 ;
        RECT 47.810 2747.020 48.990 2748.200 ;
        RECT 47.810 2568.620 48.990 2569.800 ;
        RECT 47.810 2567.020 48.990 2568.200 ;
        RECT 47.810 2388.620 48.990 2389.800 ;
        RECT 47.810 2387.020 48.990 2388.200 ;
        RECT 47.810 2208.620 48.990 2209.800 ;
        RECT 47.810 2207.020 48.990 2208.200 ;
        RECT 47.810 2028.620 48.990 2029.800 ;
        RECT 47.810 2027.020 48.990 2028.200 ;
        RECT 47.810 1848.620 48.990 1849.800 ;
        RECT 47.810 1847.020 48.990 1848.200 ;
        RECT 47.810 1668.620 48.990 1669.800 ;
        RECT 47.810 1667.020 48.990 1668.200 ;
        RECT 47.810 1488.620 48.990 1489.800 ;
        RECT 47.810 1487.020 48.990 1488.200 ;
        RECT 47.810 1308.620 48.990 1309.800 ;
        RECT 47.810 1307.020 48.990 1308.200 ;
        RECT 47.810 1128.620 48.990 1129.800 ;
        RECT 47.810 1127.020 48.990 1128.200 ;
        RECT 47.810 948.620 48.990 949.800 ;
        RECT 47.810 947.020 48.990 948.200 ;
        RECT 47.810 768.620 48.990 769.800 ;
        RECT 47.810 767.020 48.990 768.200 ;
        RECT 47.810 588.620 48.990 589.800 ;
        RECT 47.810 587.020 48.990 588.200 ;
        RECT 47.810 408.620 48.990 409.800 ;
        RECT 47.810 407.020 48.990 408.200 ;
        RECT 47.810 228.620 48.990 229.800 ;
        RECT 47.810 227.020 48.990 228.200 ;
        RECT 2970.390 3468.620 2971.570 3469.800 ;
        RECT 2970.390 3467.020 2971.570 3468.200 ;
        RECT 2970.390 3288.620 2971.570 3289.800 ;
        RECT 2970.390 3287.020 2971.570 3288.200 ;
        RECT 2970.390 3108.620 2971.570 3109.800 ;
        RECT 2970.390 3107.020 2971.570 3108.200 ;
        RECT 2970.390 2928.620 2971.570 2929.800 ;
        RECT 2970.390 2927.020 2971.570 2928.200 ;
        RECT 2970.390 2748.620 2971.570 2749.800 ;
        RECT 2970.390 2747.020 2971.570 2748.200 ;
        RECT 2970.390 2568.620 2971.570 2569.800 ;
        RECT 2970.390 2567.020 2971.570 2568.200 ;
        RECT 2970.390 2388.620 2971.570 2389.800 ;
        RECT 2970.390 2387.020 2971.570 2388.200 ;
        RECT 2970.390 2208.620 2971.570 2209.800 ;
        RECT 2970.390 2207.020 2971.570 2208.200 ;
        RECT 2970.390 2028.620 2971.570 2029.800 ;
        RECT 2970.390 2027.020 2971.570 2028.200 ;
        RECT 2970.390 1848.620 2971.570 1849.800 ;
        RECT 2970.390 1847.020 2971.570 1848.200 ;
        RECT 2970.390 1668.620 2971.570 1669.800 ;
        RECT 2970.390 1667.020 2971.570 1668.200 ;
        RECT 2970.390 1488.620 2971.570 1489.800 ;
        RECT 2970.390 1487.020 2971.570 1488.200 ;
        RECT 2970.390 1308.620 2971.570 1309.800 ;
        RECT 2970.390 1307.020 2971.570 1308.200 ;
        RECT 2970.390 1128.620 2971.570 1129.800 ;
        RECT 2970.390 1127.020 2971.570 1128.200 ;
        RECT 2970.390 948.620 2971.570 949.800 ;
        RECT 2970.390 947.020 2971.570 948.200 ;
        RECT 2970.390 768.620 2971.570 769.800 ;
        RECT 2970.390 767.020 2971.570 768.200 ;
        RECT 2970.390 588.620 2971.570 589.800 ;
        RECT 2970.390 587.020 2971.570 588.200 ;
        RECT 2970.390 408.620 2971.570 409.800 ;
        RECT 2970.390 407.020 2971.570 408.200 ;
        RECT 2970.390 228.620 2971.570 229.800 ;
        RECT 2970.390 227.020 2971.570 228.200 ;
        RECT 47.810 48.620 48.990 49.800 ;
        RECT 47.810 47.020 48.990 48.200 ;
        RECT 47.810 34.620 48.990 35.800 ;
        RECT 47.810 33.020 48.990 34.200 ;
        RECT 227.810 48.620 228.990 49.800 ;
        RECT 227.810 47.020 228.990 48.200 ;
        RECT 227.810 34.620 228.990 35.800 ;
        RECT 227.810 33.020 228.990 34.200 ;
        RECT 407.810 48.620 408.990 49.800 ;
        RECT 407.810 47.020 408.990 48.200 ;
        RECT 407.810 34.620 408.990 35.800 ;
        RECT 407.810 33.020 408.990 34.200 ;
        RECT 587.810 48.620 588.990 49.800 ;
        RECT 587.810 47.020 588.990 48.200 ;
        RECT 587.810 34.620 588.990 35.800 ;
        RECT 587.810 33.020 588.990 34.200 ;
        RECT 767.810 48.620 768.990 49.800 ;
        RECT 767.810 47.020 768.990 48.200 ;
        RECT 767.810 34.620 768.990 35.800 ;
        RECT 767.810 33.020 768.990 34.200 ;
        RECT 947.810 48.620 948.990 49.800 ;
        RECT 947.810 47.020 948.990 48.200 ;
        RECT 947.810 34.620 948.990 35.800 ;
        RECT 947.810 33.020 948.990 34.200 ;
        RECT 1127.810 48.620 1128.990 49.800 ;
        RECT 1127.810 47.020 1128.990 48.200 ;
        RECT 1127.810 34.620 1128.990 35.800 ;
        RECT 1127.810 33.020 1128.990 34.200 ;
        RECT 1307.810 48.620 1308.990 49.800 ;
        RECT 1307.810 47.020 1308.990 48.200 ;
        RECT 1307.810 34.620 1308.990 35.800 ;
        RECT 1307.810 33.020 1308.990 34.200 ;
        RECT 1487.810 48.620 1488.990 49.800 ;
        RECT 1487.810 47.020 1488.990 48.200 ;
        RECT 1487.810 34.620 1488.990 35.800 ;
        RECT 1487.810 33.020 1488.990 34.200 ;
        RECT 1667.810 48.620 1668.990 49.800 ;
        RECT 1667.810 47.020 1668.990 48.200 ;
        RECT 1667.810 34.620 1668.990 35.800 ;
        RECT 1667.810 33.020 1668.990 34.200 ;
        RECT 1847.810 48.620 1848.990 49.800 ;
        RECT 1847.810 47.020 1848.990 48.200 ;
        RECT 1847.810 34.620 1848.990 35.800 ;
        RECT 1847.810 33.020 1848.990 34.200 ;
        RECT 2027.810 48.620 2028.990 49.800 ;
        RECT 2027.810 47.020 2028.990 48.200 ;
        RECT 2027.810 34.620 2028.990 35.800 ;
        RECT 2027.810 33.020 2028.990 34.200 ;
        RECT 2207.810 48.620 2208.990 49.800 ;
        RECT 2207.810 47.020 2208.990 48.200 ;
        RECT 2207.810 34.620 2208.990 35.800 ;
        RECT 2207.810 33.020 2208.990 34.200 ;
        RECT 2387.810 48.620 2388.990 49.800 ;
        RECT 2387.810 47.020 2388.990 48.200 ;
        RECT 2387.810 34.620 2388.990 35.800 ;
        RECT 2387.810 33.020 2388.990 34.200 ;
        RECT 2567.810 48.620 2568.990 49.800 ;
        RECT 2567.810 47.020 2568.990 48.200 ;
        RECT 2567.810 34.620 2568.990 35.800 ;
        RECT 2567.810 33.020 2568.990 34.200 ;
        RECT 2747.810 48.620 2748.990 49.800 ;
        RECT 2747.810 47.020 2748.990 48.200 ;
        RECT 2747.810 34.620 2748.990 35.800 ;
        RECT 2747.810 33.020 2748.990 34.200 ;
        RECT 2927.810 48.620 2928.990 49.800 ;
        RECT 2927.810 47.020 2928.990 48.200 ;
        RECT 2927.810 34.620 2928.990 35.800 ;
        RECT 2927.810 33.020 2928.990 34.200 ;
        RECT 2970.390 48.620 2971.570 49.800 ;
        RECT 2970.390 47.020 2971.570 48.200 ;
        RECT 2970.390 34.620 2971.570 35.800 ;
        RECT 2970.390 33.020 2971.570 34.200 ;
      LAYER met5 ;
        RECT 32.900 3561.830 35.900 3561.840 ;
        RECT 46.900 3561.830 49.900 3561.840 ;
        RECT 226.900 3561.830 229.900 3561.840 ;
        RECT 406.900 3561.830 409.900 3561.840 ;
        RECT 586.900 3561.830 589.900 3561.840 ;
        RECT 766.900 3561.830 769.900 3561.840 ;
        RECT 946.900 3561.830 949.900 3561.840 ;
        RECT 1126.900 3561.830 1129.900 3561.840 ;
        RECT 1306.900 3561.830 1309.900 3561.840 ;
        RECT 1486.900 3561.830 1489.900 3561.840 ;
        RECT 1666.900 3561.830 1669.900 3561.840 ;
        RECT 1846.900 3561.830 1849.900 3561.840 ;
        RECT 2026.900 3561.830 2029.900 3561.840 ;
        RECT 2206.900 3561.830 2209.900 3561.840 ;
        RECT 2386.900 3561.830 2389.900 3561.840 ;
        RECT 2566.900 3561.830 2569.900 3561.840 ;
        RECT 2746.900 3561.830 2749.900 3561.840 ;
        RECT 2926.900 3561.830 2929.900 3561.840 ;
        RECT 2969.480 3561.830 2972.480 3561.840 ;
        RECT 32.900 3558.830 2972.480 3561.830 ;
        RECT 32.900 3558.820 35.900 3558.830 ;
        RECT 46.900 3558.820 49.900 3558.830 ;
        RECT 226.900 3558.820 229.900 3558.830 ;
        RECT 406.900 3558.820 409.900 3558.830 ;
        RECT 586.900 3558.820 589.900 3558.830 ;
        RECT 766.900 3558.820 769.900 3558.830 ;
        RECT 946.900 3558.820 949.900 3558.830 ;
        RECT 1126.900 3558.820 1129.900 3558.830 ;
        RECT 1306.900 3558.820 1309.900 3558.830 ;
        RECT 1486.900 3558.820 1489.900 3558.830 ;
        RECT 1666.900 3558.820 1669.900 3558.830 ;
        RECT 1846.900 3558.820 1849.900 3558.830 ;
        RECT 2026.900 3558.820 2029.900 3558.830 ;
        RECT 2206.900 3558.820 2209.900 3558.830 ;
        RECT 2386.900 3558.820 2389.900 3558.830 ;
        RECT 2566.900 3558.820 2569.900 3558.830 ;
        RECT 2746.900 3558.820 2749.900 3558.830 ;
        RECT 2926.900 3558.820 2929.900 3558.830 ;
        RECT 2969.480 3558.820 2972.480 3558.830 ;
        RECT 32.900 3469.910 35.900 3469.920 ;
        RECT 46.900 3469.910 49.900 3469.920 ;
        RECT 2969.480 3469.910 2972.480 3469.920 ;
        RECT 28.200 3466.910 54.000 3469.910 ;
        RECT 2951.380 3466.910 2977.180 3469.910 ;
        RECT 32.900 3466.900 35.900 3466.910 ;
        RECT 46.900 3466.900 49.900 3466.910 ;
        RECT 2969.480 3466.900 2972.480 3466.910 ;
        RECT 32.900 3289.910 35.900 3289.920 ;
        RECT 46.900 3289.910 49.900 3289.920 ;
        RECT 2969.480 3289.910 2972.480 3289.920 ;
        RECT 28.200 3286.910 54.000 3289.910 ;
        RECT 2951.380 3286.910 2977.180 3289.910 ;
        RECT 32.900 3286.900 35.900 3286.910 ;
        RECT 46.900 3286.900 49.900 3286.910 ;
        RECT 2969.480 3286.900 2972.480 3286.910 ;
        RECT 32.900 3109.910 35.900 3109.920 ;
        RECT 46.900 3109.910 49.900 3109.920 ;
        RECT 2969.480 3109.910 2972.480 3109.920 ;
        RECT 28.200 3106.910 54.000 3109.910 ;
        RECT 2951.380 3106.910 2977.180 3109.910 ;
        RECT 32.900 3106.900 35.900 3106.910 ;
        RECT 46.900 3106.900 49.900 3106.910 ;
        RECT 2969.480 3106.900 2972.480 3106.910 ;
        RECT 32.900 2929.910 35.900 2929.920 ;
        RECT 46.900 2929.910 49.900 2929.920 ;
        RECT 2969.480 2929.910 2972.480 2929.920 ;
        RECT 28.200 2926.910 54.000 2929.910 ;
        RECT 2951.380 2926.910 2977.180 2929.910 ;
        RECT 32.900 2926.900 35.900 2926.910 ;
        RECT 46.900 2926.900 49.900 2926.910 ;
        RECT 2969.480 2926.900 2972.480 2926.910 ;
        RECT 32.900 2749.910 35.900 2749.920 ;
        RECT 46.900 2749.910 49.900 2749.920 ;
        RECT 2969.480 2749.910 2972.480 2749.920 ;
        RECT 28.200 2746.910 54.000 2749.910 ;
        RECT 2951.380 2746.910 2977.180 2749.910 ;
        RECT 32.900 2746.900 35.900 2746.910 ;
        RECT 46.900 2746.900 49.900 2746.910 ;
        RECT 2969.480 2746.900 2972.480 2746.910 ;
        RECT 32.900 2569.910 35.900 2569.920 ;
        RECT 46.900 2569.910 49.900 2569.920 ;
        RECT 2969.480 2569.910 2972.480 2569.920 ;
        RECT 28.200 2566.910 54.000 2569.910 ;
        RECT 2951.380 2566.910 2977.180 2569.910 ;
        RECT 32.900 2566.900 35.900 2566.910 ;
        RECT 46.900 2566.900 49.900 2566.910 ;
        RECT 2969.480 2566.900 2972.480 2566.910 ;
        RECT 32.900 2389.910 35.900 2389.920 ;
        RECT 46.900 2389.910 49.900 2389.920 ;
        RECT 2969.480 2389.910 2972.480 2389.920 ;
        RECT 28.200 2386.910 54.000 2389.910 ;
        RECT 2951.380 2386.910 2977.180 2389.910 ;
        RECT 32.900 2386.900 35.900 2386.910 ;
        RECT 46.900 2386.900 49.900 2386.910 ;
        RECT 2969.480 2386.900 2972.480 2386.910 ;
        RECT 32.900 2209.910 35.900 2209.920 ;
        RECT 46.900 2209.910 49.900 2209.920 ;
        RECT 2969.480 2209.910 2972.480 2209.920 ;
        RECT 28.200 2206.910 54.000 2209.910 ;
        RECT 2951.380 2206.910 2977.180 2209.910 ;
        RECT 32.900 2206.900 35.900 2206.910 ;
        RECT 46.900 2206.900 49.900 2206.910 ;
        RECT 2969.480 2206.900 2972.480 2206.910 ;
        RECT 32.900 2029.910 35.900 2029.920 ;
        RECT 46.900 2029.910 49.900 2029.920 ;
        RECT 2969.480 2029.910 2972.480 2029.920 ;
        RECT 28.200 2026.910 54.000 2029.910 ;
        RECT 2951.380 2026.910 2977.180 2029.910 ;
        RECT 32.900 2026.900 35.900 2026.910 ;
        RECT 46.900 2026.900 49.900 2026.910 ;
        RECT 2969.480 2026.900 2972.480 2026.910 ;
        RECT 32.900 1849.910 35.900 1849.920 ;
        RECT 46.900 1849.910 49.900 1849.920 ;
        RECT 2969.480 1849.910 2972.480 1849.920 ;
        RECT 28.200 1846.910 54.000 1849.910 ;
        RECT 2951.380 1846.910 2977.180 1849.910 ;
        RECT 32.900 1846.900 35.900 1846.910 ;
        RECT 46.900 1846.900 49.900 1846.910 ;
        RECT 2969.480 1846.900 2972.480 1846.910 ;
        RECT 32.900 1669.910 35.900 1669.920 ;
        RECT 46.900 1669.910 49.900 1669.920 ;
        RECT 2969.480 1669.910 2972.480 1669.920 ;
        RECT 28.200 1666.910 54.000 1669.910 ;
        RECT 2951.380 1666.910 2977.180 1669.910 ;
        RECT 32.900 1666.900 35.900 1666.910 ;
        RECT 46.900 1666.900 49.900 1666.910 ;
        RECT 2969.480 1666.900 2972.480 1666.910 ;
        RECT 32.900 1489.910 35.900 1489.920 ;
        RECT 46.900 1489.910 49.900 1489.920 ;
        RECT 2969.480 1489.910 2972.480 1489.920 ;
        RECT 28.200 1486.910 54.000 1489.910 ;
        RECT 2951.380 1486.910 2977.180 1489.910 ;
        RECT 32.900 1486.900 35.900 1486.910 ;
        RECT 46.900 1486.900 49.900 1486.910 ;
        RECT 2969.480 1486.900 2972.480 1486.910 ;
        RECT 32.900 1309.910 35.900 1309.920 ;
        RECT 46.900 1309.910 49.900 1309.920 ;
        RECT 2969.480 1309.910 2972.480 1309.920 ;
        RECT 28.200 1306.910 54.000 1309.910 ;
        RECT 2951.380 1306.910 2977.180 1309.910 ;
        RECT 32.900 1306.900 35.900 1306.910 ;
        RECT 46.900 1306.900 49.900 1306.910 ;
        RECT 2969.480 1306.900 2972.480 1306.910 ;
        RECT 32.900 1129.910 35.900 1129.920 ;
        RECT 46.900 1129.910 49.900 1129.920 ;
        RECT 2969.480 1129.910 2972.480 1129.920 ;
        RECT 28.200 1126.910 54.000 1129.910 ;
        RECT 2951.380 1126.910 2977.180 1129.910 ;
        RECT 32.900 1126.900 35.900 1126.910 ;
        RECT 46.900 1126.900 49.900 1126.910 ;
        RECT 2969.480 1126.900 2972.480 1126.910 ;
        RECT 32.900 949.910 35.900 949.920 ;
        RECT 46.900 949.910 49.900 949.920 ;
        RECT 2969.480 949.910 2972.480 949.920 ;
        RECT 28.200 946.910 54.000 949.910 ;
        RECT 2951.380 946.910 2977.180 949.910 ;
        RECT 32.900 946.900 35.900 946.910 ;
        RECT 46.900 946.900 49.900 946.910 ;
        RECT 2969.480 946.900 2972.480 946.910 ;
        RECT 32.900 769.910 35.900 769.920 ;
        RECT 46.900 769.910 49.900 769.920 ;
        RECT 2969.480 769.910 2972.480 769.920 ;
        RECT 28.200 766.910 54.000 769.910 ;
        RECT 2951.380 766.910 2977.180 769.910 ;
        RECT 32.900 766.900 35.900 766.910 ;
        RECT 46.900 766.900 49.900 766.910 ;
        RECT 2969.480 766.900 2972.480 766.910 ;
        RECT 32.900 589.910 35.900 589.920 ;
        RECT 46.900 589.910 49.900 589.920 ;
        RECT 2969.480 589.910 2972.480 589.920 ;
        RECT 28.200 586.910 54.000 589.910 ;
        RECT 2951.380 586.910 2977.180 589.910 ;
        RECT 32.900 586.900 35.900 586.910 ;
        RECT 46.900 586.900 49.900 586.910 ;
        RECT 2969.480 586.900 2972.480 586.910 ;
        RECT 32.900 409.910 35.900 409.920 ;
        RECT 46.900 409.910 49.900 409.920 ;
        RECT 2969.480 409.910 2972.480 409.920 ;
        RECT 28.200 406.910 54.000 409.910 ;
        RECT 2951.380 406.910 2977.180 409.910 ;
        RECT 32.900 406.900 35.900 406.910 ;
        RECT 46.900 406.900 49.900 406.910 ;
        RECT 2969.480 406.900 2972.480 406.910 ;
        RECT 32.900 229.910 35.900 229.920 ;
        RECT 46.900 229.910 49.900 229.920 ;
        RECT 2969.480 229.910 2972.480 229.920 ;
        RECT 28.200 226.910 54.000 229.910 ;
        RECT 2951.380 226.910 2977.180 229.910 ;
        RECT 32.900 226.900 35.900 226.910 ;
        RECT 46.900 226.900 49.900 226.910 ;
        RECT 2969.480 226.900 2972.480 226.910 ;
        RECT 32.900 49.910 35.900 49.920 ;
        RECT 46.900 49.910 49.900 49.920 ;
        RECT 226.900 49.910 229.900 49.920 ;
        RECT 406.900 49.910 409.900 49.920 ;
        RECT 586.900 49.910 589.900 49.920 ;
        RECT 766.900 49.910 769.900 49.920 ;
        RECT 946.900 49.910 949.900 49.920 ;
        RECT 1126.900 49.910 1129.900 49.920 ;
        RECT 1306.900 49.910 1309.900 49.920 ;
        RECT 1486.900 49.910 1489.900 49.920 ;
        RECT 1666.900 49.910 1669.900 49.920 ;
        RECT 1846.900 49.910 1849.900 49.920 ;
        RECT 2026.900 49.910 2029.900 49.920 ;
        RECT 2206.900 49.910 2209.900 49.920 ;
        RECT 2386.900 49.910 2389.900 49.920 ;
        RECT 2566.900 49.910 2569.900 49.920 ;
        RECT 2746.900 49.910 2749.900 49.920 ;
        RECT 2926.900 49.910 2929.900 49.920 ;
        RECT 2969.480 49.910 2972.480 49.920 ;
        RECT 28.200 46.910 2977.180 49.910 ;
        RECT 32.900 46.900 35.900 46.910 ;
        RECT 46.900 46.900 49.900 46.910 ;
        RECT 226.900 46.900 229.900 46.910 ;
        RECT 406.900 46.900 409.900 46.910 ;
        RECT 586.900 46.900 589.900 46.910 ;
        RECT 766.900 46.900 769.900 46.910 ;
        RECT 946.900 46.900 949.900 46.910 ;
        RECT 1126.900 46.900 1129.900 46.910 ;
        RECT 1306.900 46.900 1309.900 46.910 ;
        RECT 1486.900 46.900 1489.900 46.910 ;
        RECT 1666.900 46.900 1669.900 46.910 ;
        RECT 1846.900 46.900 1849.900 46.910 ;
        RECT 2026.900 46.900 2029.900 46.910 ;
        RECT 2206.900 46.900 2209.900 46.910 ;
        RECT 2386.900 46.900 2389.900 46.910 ;
        RECT 2566.900 46.900 2569.900 46.910 ;
        RECT 2746.900 46.900 2749.900 46.910 ;
        RECT 2926.900 46.900 2929.900 46.910 ;
        RECT 2969.480 46.900 2972.480 46.910 ;
        RECT 32.900 35.910 35.900 35.920 ;
        RECT 46.900 35.910 49.900 35.920 ;
        RECT 226.900 35.910 229.900 35.920 ;
        RECT 406.900 35.910 409.900 35.920 ;
        RECT 586.900 35.910 589.900 35.920 ;
        RECT 766.900 35.910 769.900 35.920 ;
        RECT 946.900 35.910 949.900 35.920 ;
        RECT 1126.900 35.910 1129.900 35.920 ;
        RECT 1306.900 35.910 1309.900 35.920 ;
        RECT 1486.900 35.910 1489.900 35.920 ;
        RECT 1666.900 35.910 1669.900 35.920 ;
        RECT 1846.900 35.910 1849.900 35.920 ;
        RECT 2026.900 35.910 2029.900 35.920 ;
        RECT 2206.900 35.910 2209.900 35.920 ;
        RECT 2386.900 35.910 2389.900 35.920 ;
        RECT 2566.900 35.910 2569.900 35.920 ;
        RECT 2746.900 35.910 2749.900 35.920 ;
        RECT 2926.900 35.910 2929.900 35.920 ;
        RECT 2969.480 35.910 2972.480 35.920 ;
        RECT 32.900 32.910 2972.480 35.910 ;
        RECT 32.900 32.900 35.900 32.910 ;
        RECT 46.900 32.900 49.900 32.910 ;
        RECT 226.900 32.900 229.900 32.910 ;
        RECT 406.900 32.900 409.900 32.910 ;
        RECT 586.900 32.900 589.900 32.910 ;
        RECT 766.900 32.900 769.900 32.910 ;
        RECT 946.900 32.900 949.900 32.910 ;
        RECT 1126.900 32.900 1129.900 32.910 ;
        RECT 1306.900 32.900 1309.900 32.910 ;
        RECT 1486.900 32.900 1489.900 32.910 ;
        RECT 1666.900 32.900 1669.900 32.910 ;
        RECT 1846.900 32.900 1849.900 32.910 ;
        RECT 2026.900 32.900 2029.900 32.910 ;
        RECT 2206.900 32.900 2209.900 32.910 ;
        RECT 2386.900 32.900 2389.900 32.910 ;
        RECT 2566.900 32.900 2569.900 32.910 ;
        RECT 2746.900 32.900 2749.900 32.910 ;
        RECT 2926.900 32.900 2929.900 32.910 ;
        RECT 2969.480 32.900 2972.480 32.910 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.200 28.210 31.200 3566.530 ;
        RECT 136.900 3540.740 139.900 3566.530 ;
        RECT 316.900 3540.740 319.900 3566.530 ;
        RECT 496.900 3540.740 499.900 3566.530 ;
        RECT 676.900 3540.740 679.900 3566.530 ;
        RECT 856.900 3540.740 859.900 3566.530 ;
        RECT 1036.900 3540.740 1039.900 3566.530 ;
        RECT 1216.900 3540.740 1219.900 3566.530 ;
        RECT 1396.900 3540.740 1399.900 3566.530 ;
        RECT 1576.900 3540.740 1579.900 3566.530 ;
        RECT 1756.900 3540.740 1759.900 3566.530 ;
        RECT 1936.900 3540.740 1939.900 3566.530 ;
        RECT 2116.900 3540.740 2119.900 3566.530 ;
        RECT 2296.900 3540.740 2299.900 3566.530 ;
        RECT 2476.900 3540.740 2479.900 3566.530 ;
        RECT 2656.900 3540.740 2659.900 3566.530 ;
        RECT 2836.900 3540.740 2839.900 3566.530 ;
        RECT 136.900 28.210 139.900 54.000 ;
        RECT 316.900 28.210 319.900 54.000 ;
        RECT 496.900 28.210 499.900 54.000 ;
        RECT 676.900 28.210 679.900 54.000 ;
        RECT 856.900 28.210 859.900 54.000 ;
        RECT 1036.900 28.210 1039.900 54.000 ;
        RECT 1216.900 28.210 1219.900 54.000 ;
        RECT 1396.900 28.210 1399.900 54.000 ;
        RECT 1576.900 28.210 1579.900 54.000 ;
        RECT 1756.900 28.210 1759.900 54.000 ;
        RECT 1936.900 28.210 1939.900 54.000 ;
        RECT 2116.900 28.210 2119.900 54.000 ;
        RECT 2296.900 28.210 2299.900 54.000 ;
        RECT 2476.900 28.210 2479.900 54.000 ;
        RECT 2656.900 28.210 2659.900 54.000 ;
        RECT 2836.900 28.210 2839.900 54.000 ;
        RECT 2974.180 28.210 2977.180 3566.530 ;
      LAYER M4M5_PR_C ;
        RECT 29.110 3565.240 30.290 3566.420 ;
        RECT 29.110 3563.640 30.290 3564.820 ;
        RECT 137.810 3565.240 138.990 3566.420 ;
        RECT 137.810 3563.640 138.990 3564.820 ;
        RECT 317.810 3565.240 318.990 3566.420 ;
        RECT 317.810 3563.640 318.990 3564.820 ;
        RECT 497.810 3565.240 498.990 3566.420 ;
        RECT 497.810 3563.640 498.990 3564.820 ;
        RECT 677.810 3565.240 678.990 3566.420 ;
        RECT 677.810 3563.640 678.990 3564.820 ;
        RECT 857.810 3565.240 858.990 3566.420 ;
        RECT 857.810 3563.640 858.990 3564.820 ;
        RECT 1037.810 3565.240 1038.990 3566.420 ;
        RECT 1037.810 3563.640 1038.990 3564.820 ;
        RECT 1217.810 3565.240 1218.990 3566.420 ;
        RECT 1217.810 3563.640 1218.990 3564.820 ;
        RECT 1397.810 3565.240 1398.990 3566.420 ;
        RECT 1397.810 3563.640 1398.990 3564.820 ;
        RECT 1577.810 3565.240 1578.990 3566.420 ;
        RECT 1577.810 3563.640 1578.990 3564.820 ;
        RECT 1757.810 3565.240 1758.990 3566.420 ;
        RECT 1757.810 3563.640 1758.990 3564.820 ;
        RECT 1937.810 3565.240 1938.990 3566.420 ;
        RECT 1937.810 3563.640 1938.990 3564.820 ;
        RECT 2117.810 3565.240 2118.990 3566.420 ;
        RECT 2117.810 3563.640 2118.990 3564.820 ;
        RECT 2297.810 3565.240 2298.990 3566.420 ;
        RECT 2297.810 3563.640 2298.990 3564.820 ;
        RECT 2477.810 3565.240 2478.990 3566.420 ;
        RECT 2477.810 3563.640 2478.990 3564.820 ;
        RECT 2657.810 3565.240 2658.990 3566.420 ;
        RECT 2657.810 3563.640 2658.990 3564.820 ;
        RECT 2837.810 3565.240 2838.990 3566.420 ;
        RECT 2837.810 3563.640 2838.990 3564.820 ;
        RECT 2975.090 3565.240 2976.270 3566.420 ;
        RECT 2975.090 3563.640 2976.270 3564.820 ;
        RECT 29.110 3378.620 30.290 3379.800 ;
        RECT 29.110 3377.020 30.290 3378.200 ;
        RECT 29.110 3198.620 30.290 3199.800 ;
        RECT 29.110 3197.020 30.290 3198.200 ;
        RECT 29.110 3018.620 30.290 3019.800 ;
        RECT 29.110 3017.020 30.290 3018.200 ;
        RECT 29.110 2838.620 30.290 2839.800 ;
        RECT 29.110 2837.020 30.290 2838.200 ;
        RECT 29.110 2658.620 30.290 2659.800 ;
        RECT 29.110 2657.020 30.290 2658.200 ;
        RECT 29.110 2478.620 30.290 2479.800 ;
        RECT 29.110 2477.020 30.290 2478.200 ;
        RECT 29.110 2298.620 30.290 2299.800 ;
        RECT 29.110 2297.020 30.290 2298.200 ;
        RECT 29.110 2118.620 30.290 2119.800 ;
        RECT 29.110 2117.020 30.290 2118.200 ;
        RECT 29.110 1938.620 30.290 1939.800 ;
        RECT 29.110 1937.020 30.290 1938.200 ;
        RECT 29.110 1758.620 30.290 1759.800 ;
        RECT 29.110 1757.020 30.290 1758.200 ;
        RECT 29.110 1578.620 30.290 1579.800 ;
        RECT 29.110 1577.020 30.290 1578.200 ;
        RECT 29.110 1398.620 30.290 1399.800 ;
        RECT 29.110 1397.020 30.290 1398.200 ;
        RECT 29.110 1218.620 30.290 1219.800 ;
        RECT 29.110 1217.020 30.290 1218.200 ;
        RECT 29.110 1038.620 30.290 1039.800 ;
        RECT 29.110 1037.020 30.290 1038.200 ;
        RECT 29.110 858.620 30.290 859.800 ;
        RECT 29.110 857.020 30.290 858.200 ;
        RECT 29.110 678.620 30.290 679.800 ;
        RECT 29.110 677.020 30.290 678.200 ;
        RECT 29.110 498.620 30.290 499.800 ;
        RECT 29.110 497.020 30.290 498.200 ;
        RECT 29.110 318.620 30.290 319.800 ;
        RECT 29.110 317.020 30.290 318.200 ;
        RECT 29.110 138.620 30.290 139.800 ;
        RECT 29.110 137.020 30.290 138.200 ;
        RECT 2975.090 3378.620 2976.270 3379.800 ;
        RECT 2975.090 3377.020 2976.270 3378.200 ;
        RECT 2975.090 3198.620 2976.270 3199.800 ;
        RECT 2975.090 3197.020 2976.270 3198.200 ;
        RECT 2975.090 3018.620 2976.270 3019.800 ;
        RECT 2975.090 3017.020 2976.270 3018.200 ;
        RECT 2975.090 2838.620 2976.270 2839.800 ;
        RECT 2975.090 2837.020 2976.270 2838.200 ;
        RECT 2975.090 2658.620 2976.270 2659.800 ;
        RECT 2975.090 2657.020 2976.270 2658.200 ;
        RECT 2975.090 2478.620 2976.270 2479.800 ;
        RECT 2975.090 2477.020 2976.270 2478.200 ;
        RECT 2975.090 2298.620 2976.270 2299.800 ;
        RECT 2975.090 2297.020 2976.270 2298.200 ;
        RECT 2975.090 2118.620 2976.270 2119.800 ;
        RECT 2975.090 2117.020 2976.270 2118.200 ;
        RECT 2975.090 1938.620 2976.270 1939.800 ;
        RECT 2975.090 1937.020 2976.270 1938.200 ;
        RECT 2975.090 1758.620 2976.270 1759.800 ;
        RECT 2975.090 1757.020 2976.270 1758.200 ;
        RECT 2975.090 1578.620 2976.270 1579.800 ;
        RECT 2975.090 1577.020 2976.270 1578.200 ;
        RECT 2975.090 1398.620 2976.270 1399.800 ;
        RECT 2975.090 1397.020 2976.270 1398.200 ;
        RECT 2975.090 1218.620 2976.270 1219.800 ;
        RECT 2975.090 1217.020 2976.270 1218.200 ;
        RECT 2975.090 1038.620 2976.270 1039.800 ;
        RECT 2975.090 1037.020 2976.270 1038.200 ;
        RECT 2975.090 858.620 2976.270 859.800 ;
        RECT 2975.090 857.020 2976.270 858.200 ;
        RECT 2975.090 678.620 2976.270 679.800 ;
        RECT 2975.090 677.020 2976.270 678.200 ;
        RECT 2975.090 498.620 2976.270 499.800 ;
        RECT 2975.090 497.020 2976.270 498.200 ;
        RECT 2975.090 318.620 2976.270 319.800 ;
        RECT 2975.090 317.020 2976.270 318.200 ;
        RECT 2975.090 138.620 2976.270 139.800 ;
        RECT 2975.090 137.020 2976.270 138.200 ;
        RECT 29.110 29.920 30.290 31.100 ;
        RECT 29.110 28.320 30.290 29.500 ;
        RECT 137.810 29.920 138.990 31.100 ;
        RECT 137.810 28.320 138.990 29.500 ;
        RECT 317.810 29.920 318.990 31.100 ;
        RECT 317.810 28.320 318.990 29.500 ;
        RECT 497.810 29.920 498.990 31.100 ;
        RECT 497.810 28.320 498.990 29.500 ;
        RECT 677.810 29.920 678.990 31.100 ;
        RECT 677.810 28.320 678.990 29.500 ;
        RECT 857.810 29.920 858.990 31.100 ;
        RECT 857.810 28.320 858.990 29.500 ;
        RECT 1037.810 29.920 1038.990 31.100 ;
        RECT 1037.810 28.320 1038.990 29.500 ;
        RECT 1217.810 29.920 1218.990 31.100 ;
        RECT 1217.810 28.320 1218.990 29.500 ;
        RECT 1397.810 29.920 1398.990 31.100 ;
        RECT 1397.810 28.320 1398.990 29.500 ;
        RECT 1577.810 29.920 1578.990 31.100 ;
        RECT 1577.810 28.320 1578.990 29.500 ;
        RECT 1757.810 29.920 1758.990 31.100 ;
        RECT 1757.810 28.320 1758.990 29.500 ;
        RECT 1937.810 29.920 1938.990 31.100 ;
        RECT 1937.810 28.320 1938.990 29.500 ;
        RECT 2117.810 29.920 2118.990 31.100 ;
        RECT 2117.810 28.320 2118.990 29.500 ;
        RECT 2297.810 29.920 2298.990 31.100 ;
        RECT 2297.810 28.320 2298.990 29.500 ;
        RECT 2477.810 29.920 2478.990 31.100 ;
        RECT 2477.810 28.320 2478.990 29.500 ;
        RECT 2657.810 29.920 2658.990 31.100 ;
        RECT 2657.810 28.320 2658.990 29.500 ;
        RECT 2837.810 29.920 2838.990 31.100 ;
        RECT 2837.810 28.320 2838.990 29.500 ;
        RECT 2975.090 29.920 2976.270 31.100 ;
        RECT 2975.090 28.320 2976.270 29.500 ;
      LAYER met5 ;
        RECT 28.200 3566.530 31.200 3566.540 ;
        RECT 136.900 3566.530 139.900 3566.540 ;
        RECT 316.900 3566.530 319.900 3566.540 ;
        RECT 496.900 3566.530 499.900 3566.540 ;
        RECT 676.900 3566.530 679.900 3566.540 ;
        RECT 856.900 3566.530 859.900 3566.540 ;
        RECT 1036.900 3566.530 1039.900 3566.540 ;
        RECT 1216.900 3566.530 1219.900 3566.540 ;
        RECT 1396.900 3566.530 1399.900 3566.540 ;
        RECT 1576.900 3566.530 1579.900 3566.540 ;
        RECT 1756.900 3566.530 1759.900 3566.540 ;
        RECT 1936.900 3566.530 1939.900 3566.540 ;
        RECT 2116.900 3566.530 2119.900 3566.540 ;
        RECT 2296.900 3566.530 2299.900 3566.540 ;
        RECT 2476.900 3566.530 2479.900 3566.540 ;
        RECT 2656.900 3566.530 2659.900 3566.540 ;
        RECT 2836.900 3566.530 2839.900 3566.540 ;
        RECT 2974.180 3566.530 2977.180 3566.540 ;
        RECT 28.200 3563.530 2977.180 3566.530 ;
        RECT 28.200 3563.520 31.200 3563.530 ;
        RECT 136.900 3563.520 139.900 3563.530 ;
        RECT 316.900 3563.520 319.900 3563.530 ;
        RECT 496.900 3563.520 499.900 3563.530 ;
        RECT 676.900 3563.520 679.900 3563.530 ;
        RECT 856.900 3563.520 859.900 3563.530 ;
        RECT 1036.900 3563.520 1039.900 3563.530 ;
        RECT 1216.900 3563.520 1219.900 3563.530 ;
        RECT 1396.900 3563.520 1399.900 3563.530 ;
        RECT 1576.900 3563.520 1579.900 3563.530 ;
        RECT 1756.900 3563.520 1759.900 3563.530 ;
        RECT 1936.900 3563.520 1939.900 3563.530 ;
        RECT 2116.900 3563.520 2119.900 3563.530 ;
        RECT 2296.900 3563.520 2299.900 3563.530 ;
        RECT 2476.900 3563.520 2479.900 3563.530 ;
        RECT 2656.900 3563.520 2659.900 3563.530 ;
        RECT 2836.900 3563.520 2839.900 3563.530 ;
        RECT 2974.180 3563.520 2977.180 3563.530 ;
        RECT 28.200 3379.910 31.200 3379.920 ;
        RECT 2974.180 3379.910 2977.180 3379.920 ;
        RECT 28.200 3376.910 54.000 3379.910 ;
        RECT 2951.380 3376.910 2977.180 3379.910 ;
        RECT 28.200 3376.900 31.200 3376.910 ;
        RECT 2974.180 3376.900 2977.180 3376.910 ;
        RECT 28.200 3199.910 31.200 3199.920 ;
        RECT 2974.180 3199.910 2977.180 3199.920 ;
        RECT 28.200 3196.910 54.000 3199.910 ;
        RECT 2951.380 3196.910 2977.180 3199.910 ;
        RECT 28.200 3196.900 31.200 3196.910 ;
        RECT 2974.180 3196.900 2977.180 3196.910 ;
        RECT 28.200 3019.910 31.200 3019.920 ;
        RECT 2974.180 3019.910 2977.180 3019.920 ;
        RECT 28.200 3016.910 54.000 3019.910 ;
        RECT 2951.380 3016.910 2977.180 3019.910 ;
        RECT 28.200 3016.900 31.200 3016.910 ;
        RECT 2974.180 3016.900 2977.180 3016.910 ;
        RECT 28.200 2839.910 31.200 2839.920 ;
        RECT 2974.180 2839.910 2977.180 2839.920 ;
        RECT 28.200 2836.910 54.000 2839.910 ;
        RECT 2951.380 2836.910 2977.180 2839.910 ;
        RECT 28.200 2836.900 31.200 2836.910 ;
        RECT 2974.180 2836.900 2977.180 2836.910 ;
        RECT 28.200 2659.910 31.200 2659.920 ;
        RECT 2974.180 2659.910 2977.180 2659.920 ;
        RECT 28.200 2656.910 54.000 2659.910 ;
        RECT 2951.380 2656.910 2977.180 2659.910 ;
        RECT 28.200 2656.900 31.200 2656.910 ;
        RECT 2974.180 2656.900 2977.180 2656.910 ;
        RECT 28.200 2479.910 31.200 2479.920 ;
        RECT 2974.180 2479.910 2977.180 2479.920 ;
        RECT 28.200 2476.910 54.000 2479.910 ;
        RECT 2951.380 2476.910 2977.180 2479.910 ;
        RECT 28.200 2476.900 31.200 2476.910 ;
        RECT 2974.180 2476.900 2977.180 2476.910 ;
        RECT 28.200 2299.910 31.200 2299.920 ;
        RECT 2974.180 2299.910 2977.180 2299.920 ;
        RECT 28.200 2296.910 54.000 2299.910 ;
        RECT 2951.380 2296.910 2977.180 2299.910 ;
        RECT 28.200 2296.900 31.200 2296.910 ;
        RECT 2974.180 2296.900 2977.180 2296.910 ;
        RECT 28.200 2119.910 31.200 2119.920 ;
        RECT 2974.180 2119.910 2977.180 2119.920 ;
        RECT 28.200 2116.910 54.000 2119.910 ;
        RECT 2951.380 2116.910 2977.180 2119.910 ;
        RECT 28.200 2116.900 31.200 2116.910 ;
        RECT 2974.180 2116.900 2977.180 2116.910 ;
        RECT 28.200 1939.910 31.200 1939.920 ;
        RECT 2974.180 1939.910 2977.180 1939.920 ;
        RECT 28.200 1936.910 54.000 1939.910 ;
        RECT 2951.380 1936.910 2977.180 1939.910 ;
        RECT 28.200 1936.900 31.200 1936.910 ;
        RECT 2974.180 1936.900 2977.180 1936.910 ;
        RECT 28.200 1759.910 31.200 1759.920 ;
        RECT 2974.180 1759.910 2977.180 1759.920 ;
        RECT 28.200 1756.910 54.000 1759.910 ;
        RECT 2951.380 1756.910 2977.180 1759.910 ;
        RECT 28.200 1756.900 31.200 1756.910 ;
        RECT 2974.180 1756.900 2977.180 1756.910 ;
        RECT 28.200 1579.910 31.200 1579.920 ;
        RECT 2974.180 1579.910 2977.180 1579.920 ;
        RECT 28.200 1576.910 54.000 1579.910 ;
        RECT 2951.380 1576.910 2977.180 1579.910 ;
        RECT 28.200 1576.900 31.200 1576.910 ;
        RECT 2974.180 1576.900 2977.180 1576.910 ;
        RECT 28.200 1399.910 31.200 1399.920 ;
        RECT 2974.180 1399.910 2977.180 1399.920 ;
        RECT 28.200 1396.910 54.000 1399.910 ;
        RECT 2951.380 1396.910 2977.180 1399.910 ;
        RECT 28.200 1396.900 31.200 1396.910 ;
        RECT 2974.180 1396.900 2977.180 1396.910 ;
        RECT 28.200 1219.910 31.200 1219.920 ;
        RECT 2974.180 1219.910 2977.180 1219.920 ;
        RECT 28.200 1216.910 54.000 1219.910 ;
        RECT 2951.380 1216.910 2977.180 1219.910 ;
        RECT 28.200 1216.900 31.200 1216.910 ;
        RECT 2974.180 1216.900 2977.180 1216.910 ;
        RECT 28.200 1039.910 31.200 1039.920 ;
        RECT 2974.180 1039.910 2977.180 1039.920 ;
        RECT 28.200 1036.910 54.000 1039.910 ;
        RECT 2951.380 1036.910 2977.180 1039.910 ;
        RECT 28.200 1036.900 31.200 1036.910 ;
        RECT 2974.180 1036.900 2977.180 1036.910 ;
        RECT 28.200 859.910 31.200 859.920 ;
        RECT 2974.180 859.910 2977.180 859.920 ;
        RECT 28.200 856.910 54.000 859.910 ;
        RECT 2951.380 856.910 2977.180 859.910 ;
        RECT 28.200 856.900 31.200 856.910 ;
        RECT 2974.180 856.900 2977.180 856.910 ;
        RECT 28.200 679.910 31.200 679.920 ;
        RECT 2974.180 679.910 2977.180 679.920 ;
        RECT 28.200 676.910 54.000 679.910 ;
        RECT 2951.380 676.910 2977.180 679.910 ;
        RECT 28.200 676.900 31.200 676.910 ;
        RECT 2974.180 676.900 2977.180 676.910 ;
        RECT 28.200 499.910 31.200 499.920 ;
        RECT 2974.180 499.910 2977.180 499.920 ;
        RECT 28.200 496.910 54.000 499.910 ;
        RECT 2951.380 496.910 2977.180 499.910 ;
        RECT 28.200 496.900 31.200 496.910 ;
        RECT 2974.180 496.900 2977.180 496.910 ;
        RECT 28.200 319.910 31.200 319.920 ;
        RECT 2974.180 319.910 2977.180 319.920 ;
        RECT 28.200 316.910 54.000 319.910 ;
        RECT 2951.380 316.910 2977.180 319.910 ;
        RECT 28.200 316.900 31.200 316.910 ;
        RECT 2974.180 316.900 2977.180 316.910 ;
        RECT 28.200 139.910 31.200 139.920 ;
        RECT 2974.180 139.910 2977.180 139.920 ;
        RECT 28.200 136.910 54.000 139.910 ;
        RECT 2951.380 136.910 2977.180 139.910 ;
        RECT 28.200 136.900 31.200 136.910 ;
        RECT 2974.180 136.900 2977.180 136.910 ;
        RECT 28.200 31.210 31.200 31.220 ;
        RECT 136.900 31.210 139.900 31.220 ;
        RECT 316.900 31.210 319.900 31.220 ;
        RECT 496.900 31.210 499.900 31.220 ;
        RECT 676.900 31.210 679.900 31.220 ;
        RECT 856.900 31.210 859.900 31.220 ;
        RECT 1036.900 31.210 1039.900 31.220 ;
        RECT 1216.900 31.210 1219.900 31.220 ;
        RECT 1396.900 31.210 1399.900 31.220 ;
        RECT 1576.900 31.210 1579.900 31.220 ;
        RECT 1756.900 31.210 1759.900 31.220 ;
        RECT 1936.900 31.210 1939.900 31.220 ;
        RECT 2116.900 31.210 2119.900 31.220 ;
        RECT 2296.900 31.210 2299.900 31.220 ;
        RECT 2476.900 31.210 2479.900 31.220 ;
        RECT 2656.900 31.210 2659.900 31.220 ;
        RECT 2836.900 31.210 2839.900 31.220 ;
        RECT 2974.180 31.210 2977.180 31.220 ;
        RECT 28.200 28.210 2977.180 31.210 ;
        RECT 28.200 28.200 31.200 28.210 ;
        RECT 136.900 28.200 139.900 28.210 ;
        RECT 316.900 28.200 319.900 28.210 ;
        RECT 496.900 28.200 499.900 28.210 ;
        RECT 676.900 28.200 679.900 28.210 ;
        RECT 856.900 28.200 859.900 28.210 ;
        RECT 1036.900 28.200 1039.900 28.210 ;
        RECT 1216.900 28.200 1219.900 28.210 ;
        RECT 1396.900 28.200 1399.900 28.210 ;
        RECT 1576.900 28.200 1579.900 28.210 ;
        RECT 1756.900 28.200 1759.900 28.210 ;
        RECT 1936.900 28.200 1939.900 28.210 ;
        RECT 2116.900 28.200 2119.900 28.210 ;
        RECT 2296.900 28.200 2299.900 28.210 ;
        RECT 2476.900 28.200 2479.900 28.210 ;
        RECT 2656.900 28.200 2659.900 28.210 ;
        RECT 2836.900 28.200 2839.900 28.210 ;
        RECT 2974.180 28.200 2977.180 28.210 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 23.500 23.510 26.500 3571.230 ;
        RECT 2978.880 23.510 2981.880 3571.230 ;
      LAYER M4M5_PR_C ;
        RECT 24.410 3569.940 25.590 3571.120 ;
        RECT 24.410 3568.340 25.590 3569.520 ;
        RECT 24.410 25.220 25.590 26.400 ;
        RECT 24.410 23.620 25.590 24.800 ;
        RECT 2979.790 3569.940 2980.970 3571.120 ;
        RECT 2979.790 3568.340 2980.970 3569.520 ;
        RECT 2979.790 25.220 2980.970 26.400 ;
        RECT 2979.790 23.620 2980.970 24.800 ;
      LAYER met5 ;
        RECT 23.500 3571.230 26.500 3571.240 ;
        RECT 2978.880 3571.230 2981.880 3571.240 ;
        RECT 23.500 3568.230 2981.880 3571.230 ;
        RECT 23.500 3568.220 26.500 3568.230 ;
        RECT 2978.880 3568.220 2981.880 3568.230 ;
        RECT 23.500 26.510 26.500 26.520 ;
        RECT 2978.880 26.510 2981.880 26.520 ;
        RECT 23.500 23.510 2981.880 26.510 ;
        RECT 23.500 23.500 26.500 23.510 ;
        RECT 2978.880 23.500 2981.880 23.510 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 18.800 18.810 21.800 3575.930 ;
        RECT 2983.580 18.810 2986.580 3575.930 ;
      LAYER M4M5_PR_C ;
        RECT 19.710 3574.640 20.890 3575.820 ;
        RECT 19.710 3573.040 20.890 3574.220 ;
        RECT 19.710 20.520 20.890 21.700 ;
        RECT 19.710 18.920 20.890 20.100 ;
        RECT 2984.490 3574.640 2985.670 3575.820 ;
        RECT 2984.490 3573.040 2985.670 3574.220 ;
        RECT 2984.490 20.520 2985.670 21.700 ;
        RECT 2984.490 18.920 2985.670 20.100 ;
      LAYER met5 ;
        RECT 18.800 3575.930 21.800 3575.940 ;
        RECT 2983.580 3575.930 2986.580 3575.940 ;
        RECT 18.800 3572.930 2986.580 3575.930 ;
        RECT 18.800 3572.920 21.800 3572.930 ;
        RECT 2983.580 3572.920 2986.580 3572.930 ;
        RECT 18.800 21.810 21.800 21.820 ;
        RECT 2983.580 21.810 2986.580 21.820 ;
        RECT 18.800 18.810 2986.580 21.810 ;
        RECT 18.800 18.800 21.800 18.810 ;
        RECT 2983.580 18.800 2986.580 18.810 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 14.100 14.110 17.100 3580.630 ;
        RECT 2988.280 14.110 2991.280 3580.630 ;
      LAYER M4M5_PR_C ;
        RECT 15.010 3579.340 16.190 3580.520 ;
        RECT 15.010 3577.740 16.190 3578.920 ;
        RECT 15.010 15.820 16.190 17.000 ;
        RECT 15.010 14.220 16.190 15.400 ;
        RECT 2989.190 3579.340 2990.370 3580.520 ;
        RECT 2989.190 3577.740 2990.370 3578.920 ;
        RECT 2989.190 15.820 2990.370 17.000 ;
        RECT 2989.190 14.220 2990.370 15.400 ;
      LAYER met5 ;
        RECT 14.100 3580.630 17.100 3580.640 ;
        RECT 2988.280 3580.630 2991.280 3580.640 ;
        RECT 14.100 3577.630 2991.280 3580.630 ;
        RECT 14.100 3577.620 17.100 3577.630 ;
        RECT 2988.280 3577.620 2991.280 3577.630 ;
        RECT 14.100 17.110 17.100 17.120 ;
        RECT 2988.280 17.110 2991.280 17.120 ;
        RECT 14.100 14.110 2991.280 17.110 ;
        RECT 14.100 14.100 17.100 14.110 ;
        RECT 2988.280 14.100 2991.280 14.110 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 9.400 9.410 12.400 3585.330 ;
        RECT 2992.980 9.410 2995.980 3585.330 ;
      LAYER M4M5_PR_C ;
        RECT 10.310 3584.040 11.490 3585.220 ;
        RECT 10.310 3582.440 11.490 3583.620 ;
        RECT 10.310 11.120 11.490 12.300 ;
        RECT 10.310 9.520 11.490 10.700 ;
        RECT 2993.890 3584.040 2995.070 3585.220 ;
        RECT 2993.890 3582.440 2995.070 3583.620 ;
        RECT 2993.890 11.120 2995.070 12.300 ;
        RECT 2993.890 9.520 2995.070 10.700 ;
      LAYER met5 ;
        RECT 9.400 3585.330 12.400 3585.340 ;
        RECT 2992.980 3585.330 2995.980 3585.340 ;
        RECT 9.400 3582.330 2995.980 3585.330 ;
        RECT 9.400 3582.320 12.400 3582.330 ;
        RECT 2992.980 3582.320 2995.980 3582.330 ;
        RECT 9.400 12.410 12.400 12.420 ;
        RECT 2992.980 12.410 2995.980 12.420 ;
        RECT 9.400 9.410 2995.980 12.410 ;
        RECT 9.400 9.400 12.400 9.410 ;
        RECT 2992.980 9.400 2995.980 9.410 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 4.700 4.710 7.700 3590.030 ;
        RECT 2997.680 4.710 3000.680 3590.030 ;
      LAYER M4M5_PR_C ;
        RECT 5.610 3588.740 6.790 3589.920 ;
        RECT 5.610 3587.140 6.790 3588.320 ;
        RECT 5.610 6.420 6.790 7.600 ;
        RECT 5.610 4.820 6.790 6.000 ;
        RECT 2998.590 3588.740 2999.770 3589.920 ;
        RECT 2998.590 3587.140 2999.770 3588.320 ;
        RECT 2998.590 6.420 2999.770 7.600 ;
        RECT 2998.590 4.820 2999.770 6.000 ;
      LAYER met5 ;
        RECT 4.700 3590.030 7.700 3590.040 ;
        RECT 2997.680 3590.030 3000.680 3590.040 ;
        RECT 4.700 3587.030 3000.680 3590.030 ;
        RECT 4.700 3587.020 7.700 3587.030 ;
        RECT 2997.680 3587.020 3000.680 3587.030 ;
        RECT 4.700 7.710 7.700 7.720 ;
        RECT 2997.680 7.710 3000.680 7.720 ;
        RECT 4.700 4.710 3000.680 7.710 ;
        RECT 4.700 4.700 7.700 4.710 ;
        RECT 2997.680 4.700 3000.680 4.710 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.010 3.000 3594.730 ;
        RECT 3002.380 0.010 3005.380 3594.730 ;
      LAYER M4M5_PR_C ;
        RECT 0.910 3593.440 2.090 3594.620 ;
        RECT 0.910 3591.840 2.090 3593.020 ;
        RECT 0.910 1.720 2.090 2.900 ;
        RECT 0.910 0.120 2.090 1.300 ;
        RECT 3003.290 3593.440 3004.470 3594.620 ;
        RECT 3003.290 3591.840 3004.470 3593.020 ;
        RECT 3003.290 1.720 3004.470 2.900 ;
        RECT 3003.290 0.120 3004.470 1.300 ;
      LAYER met5 ;
        RECT 0.000 3594.730 3.000 3594.740 ;
        RECT 3002.380 3594.730 3005.380 3594.740 ;
        RECT 0.000 3591.730 3005.380 3594.730 ;
        RECT 0.000 3591.720 3.000 3591.730 ;
        RECT 3002.380 3591.720 3005.380 3591.730 ;
        RECT 0.000 3.010 3.000 3.020 ;
        RECT 3002.380 3.010 3005.380 3.020 ;
        RECT 0.000 0.010 3005.380 3.010 ;
        RECT 0.000 0.000 3.000 0.010 ;
        RECT 3002.380 0.000 3005.380 0.010 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 697.625 369.205 2441.635 3266.765 ;
      LAYER met1 ;
        RECT 54.000 54.000 2944.490 3540.740 ;
      LAYER met2 ;
        RECT 56.320 54.000 2947.690 3540.740 ;
      LAYER met3 ;
        RECT 54.000 73.065 2951.380 3539.355 ;
      LAYER met4 ;
        RECT 136.900 54.000 2929.900 3540.740 ;
      LAYER met5 ;
        RECT 54.000 136.900 2951.380 3469.920 ;
  END
END user_project_wrapper
END LIBRARY

