VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pyfive_top
  CLASS BLOCK ;
  FOREIGN pyfive_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 1748.000 BY 1360.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 13.640 1748.000 14.240 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 863.640 1748.000 864.240 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 948.640 1748.000 949.240 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 1033.640 1748.000 1034.240 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 1118.640 1748.000 1119.240 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 1203.640 1748.000 1204.240 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 1288.640 1748.000 1289.240 ;
    END
  END io_in[15]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 98.640 1748.000 99.240 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 183.640 1748.000 184.240 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 268.640 1748.000 269.240 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 353.640 1748.000 354.240 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 438.640 1748.000 439.240 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 523.640 1748.000 524.240 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 608.640 1748.000 609.240 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 693.640 1748.000 694.240 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1744.000 778.640 1748.000 779.240 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 41.520 1748.000 42.120 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 891.520 1748.000 892.120 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 976.520 1748.000 977.120 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 1061.520 1748.000 1062.120 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 1146.520 1748.000 1147.120 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 1231.520 1748.000 1232.120 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 1316.520 1748.000 1317.120 ;
    END
  END io_oeb[15]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 126.520 1748.000 127.120 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 211.520 1748.000 212.120 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 296.520 1748.000 297.120 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 381.520 1748.000 382.120 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 466.520 1748.000 467.120 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 551.520 1748.000 552.120 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 636.520 1748.000 637.120 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 721.520 1748.000 722.120 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 806.520 1748.000 807.120 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 70.080 1748.000 70.680 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 920.080 1748.000 920.680 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 1005.080 1748.000 1005.680 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 1090.080 1748.000 1090.680 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 1175.080 1748.000 1175.680 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 1260.080 1748.000 1260.680 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 1345.080 1748.000 1345.680 ;
    END
  END io_out[15]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 155.080 1748.000 155.680 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 240.080 1748.000 240.680 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 325.080 1748.000 325.680 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 410.080 1748.000 410.680 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 495.080 1748.000 495.680 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 580.080 1748.000 580.680 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 665.080 1748.000 665.680 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 750.080 1748.000 750.680 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1744.000 835.080 1748.000 835.680 ;
    END
  END io_out[9]
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1311.090 1356.000 1311.370 1360.000 ;
    END
  END one
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.880 4.000 519.480 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 634.480 4.000 635.080 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 711.320 4.000 711.920 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 750.080 4.000 750.680 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.160 4.000 788.760 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.920 4.000 827.520 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.680 4.000 866.280 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 903.760 4.000 904.360 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 942.520 4.000 943.120 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1019.360 4.000 1019.960 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1058.120 4.000 1058.720 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1096.200 4.000 1096.800 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1134.960 4.000 1135.560 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.040 4.000 1173.640 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1211.800 4.000 1212.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1250.560 4.000 1251.160 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1288.640 4.000 1289.240 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1327.400 4.000 1328.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.200 4.000 365.800 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.280 4.000 403.880 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.800 4.000 481.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 570.560 4.000 571.160 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.160 4.000 686.760 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.000 4.000 763.600 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.080 4.000 801.680 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 878.600 4.000 879.200 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.680 4.000 917.280 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 993.520 4.000 994.120 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1032.280 4.000 1032.880 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.040 4.000 1071.640 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1109.120 4.000 1109.720 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1147.880 4.000 1148.480 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1185.960 4.000 1186.560 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1224.720 4.000 1225.320 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1263.480 4.000 1264.080 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1301.560 4.000 1302.160 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1340.320 4.000 1340.920 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.960 4.000 455.560 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.720 4.000 545.320 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 698.400 4.000 699.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.160 4.000 737.760 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.920 4.000 776.520 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.000 4.000 814.600 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 852.760 4.000 853.360 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.840 4.000 891.440 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 929.600 4.000 930.200 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 968.360 4.000 968.960 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1006.440 4.000 1007.040 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1045.200 4.000 1045.800 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1083.280 4.000 1083.880 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 4.000 1122.640 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1160.800 4.000 1161.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1198.880 4.000 1199.480 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1237.640 4.000 1238.240 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.720 4.000 1276.320 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1314.480 4.000 1315.080 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1353.240 4.000 1353.840 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.520 4.000 314.120 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.960 4.000 506.560 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END wbs_we_i
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 437.090 1356.000 437.370 1360.000 ;
    END
  END zero
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 49.200 1742.480 50.800 ;
        RECT 5.520 228.200 1742.480 230.800 ;
        RECT 5.520 408.200 1742.480 410.800 ;
        RECT 5.520 588.200 1742.480 590.800 ;
        RECT 5.520 768.200 1742.480 770.800 ;
        RECT 5.520 948.200 1742.480 950.800 ;
        RECT 5.520 1128.200 1742.480 1130.800 ;
        RECT 5.520 1308.200 1742.480 1310.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 139.200 1742.480 140.800 ;
        RECT 5.520 319.200 1742.480 320.800 ;
        RECT 5.520 499.200 1742.480 500.800 ;
        RECT 5.520 679.200 1742.480 680.800 ;
        RECT 5.520 859.200 1742.480 860.800 ;
        RECT 5.520 1039.200 1742.480 1040.800 ;
        RECT 5.520 1219.200 1742.480 1220.800 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1742.480 1349.205 ;
      LAYER met1 ;
        RECT 3.750 6.500 1742.480 1349.360 ;
      LAYER met2 ;
        RECT 3.780 1355.720 436.810 1356.000 ;
        RECT 437.650 1355.720 1310.810 1356.000 ;
        RECT 1311.650 1355.720 1736.110 1356.000 ;
        RECT 3.780 6.275 1736.110 1355.720 ;
      LAYER met3 ;
        RECT 4.400 1352.840 1744.010 1353.705 ;
        RECT 4.000 1346.080 1744.010 1352.840 ;
        RECT 4.000 1344.680 1743.600 1346.080 ;
        RECT 4.000 1341.320 1744.010 1344.680 ;
        RECT 4.400 1339.920 1744.010 1341.320 ;
        RECT 4.000 1328.400 1744.010 1339.920 ;
        RECT 4.400 1327.000 1744.010 1328.400 ;
        RECT 4.000 1317.520 1744.010 1327.000 ;
        RECT 4.000 1316.120 1743.600 1317.520 ;
        RECT 4.000 1315.480 1744.010 1316.120 ;
        RECT 4.400 1314.080 1744.010 1315.480 ;
        RECT 4.000 1302.560 1744.010 1314.080 ;
        RECT 4.400 1301.160 1744.010 1302.560 ;
        RECT 4.000 1289.640 1744.010 1301.160 ;
        RECT 4.400 1288.240 1743.600 1289.640 ;
        RECT 4.000 1276.720 1744.010 1288.240 ;
        RECT 4.400 1275.320 1744.010 1276.720 ;
        RECT 4.000 1264.480 1744.010 1275.320 ;
        RECT 4.400 1263.080 1744.010 1264.480 ;
        RECT 4.000 1261.080 1744.010 1263.080 ;
        RECT 4.000 1259.680 1743.600 1261.080 ;
        RECT 4.000 1251.560 1744.010 1259.680 ;
        RECT 4.400 1250.160 1744.010 1251.560 ;
        RECT 4.000 1238.640 1744.010 1250.160 ;
        RECT 4.400 1237.240 1744.010 1238.640 ;
        RECT 4.000 1232.520 1744.010 1237.240 ;
        RECT 4.000 1231.120 1743.600 1232.520 ;
        RECT 4.000 1225.720 1744.010 1231.120 ;
        RECT 4.400 1224.320 1744.010 1225.720 ;
        RECT 4.000 1212.800 1744.010 1224.320 ;
        RECT 4.400 1211.400 1744.010 1212.800 ;
        RECT 4.000 1204.640 1744.010 1211.400 ;
        RECT 4.000 1203.240 1743.600 1204.640 ;
        RECT 4.000 1199.880 1744.010 1203.240 ;
        RECT 4.400 1198.480 1744.010 1199.880 ;
        RECT 4.000 1186.960 1744.010 1198.480 ;
        RECT 4.400 1185.560 1744.010 1186.960 ;
        RECT 4.000 1176.080 1744.010 1185.560 ;
        RECT 4.000 1174.680 1743.600 1176.080 ;
        RECT 4.000 1174.040 1744.010 1174.680 ;
        RECT 4.400 1172.640 1744.010 1174.040 ;
        RECT 4.000 1161.800 1744.010 1172.640 ;
        RECT 4.400 1160.400 1744.010 1161.800 ;
        RECT 4.000 1148.880 1744.010 1160.400 ;
        RECT 4.400 1147.520 1744.010 1148.880 ;
        RECT 4.400 1147.480 1743.600 1147.520 ;
        RECT 4.000 1146.120 1743.600 1147.480 ;
        RECT 4.000 1135.960 1744.010 1146.120 ;
        RECT 4.400 1134.560 1744.010 1135.960 ;
        RECT 4.000 1123.040 1744.010 1134.560 ;
        RECT 4.400 1121.640 1744.010 1123.040 ;
        RECT 4.000 1119.640 1744.010 1121.640 ;
        RECT 4.000 1118.240 1743.600 1119.640 ;
        RECT 4.000 1110.120 1744.010 1118.240 ;
        RECT 4.400 1108.720 1744.010 1110.120 ;
        RECT 4.000 1097.200 1744.010 1108.720 ;
        RECT 4.400 1095.800 1744.010 1097.200 ;
        RECT 4.000 1091.080 1744.010 1095.800 ;
        RECT 4.000 1089.680 1743.600 1091.080 ;
        RECT 4.000 1084.280 1744.010 1089.680 ;
        RECT 4.400 1082.880 1744.010 1084.280 ;
        RECT 4.000 1072.040 1744.010 1082.880 ;
        RECT 4.400 1070.640 1744.010 1072.040 ;
        RECT 4.000 1062.520 1744.010 1070.640 ;
        RECT 4.000 1061.120 1743.600 1062.520 ;
        RECT 4.000 1059.120 1744.010 1061.120 ;
        RECT 4.400 1057.720 1744.010 1059.120 ;
        RECT 4.000 1046.200 1744.010 1057.720 ;
        RECT 4.400 1044.800 1744.010 1046.200 ;
        RECT 4.000 1034.640 1744.010 1044.800 ;
        RECT 4.000 1033.280 1743.600 1034.640 ;
        RECT 4.400 1033.240 1743.600 1033.280 ;
        RECT 4.400 1031.880 1744.010 1033.240 ;
        RECT 4.000 1020.360 1744.010 1031.880 ;
        RECT 4.400 1018.960 1744.010 1020.360 ;
        RECT 4.000 1007.440 1744.010 1018.960 ;
        RECT 4.400 1006.080 1744.010 1007.440 ;
        RECT 4.400 1006.040 1743.600 1006.080 ;
        RECT 4.000 1004.680 1743.600 1006.040 ;
        RECT 4.000 994.520 1744.010 1004.680 ;
        RECT 4.400 993.120 1744.010 994.520 ;
        RECT 4.000 981.600 1744.010 993.120 ;
        RECT 4.400 980.200 1744.010 981.600 ;
        RECT 4.000 977.520 1744.010 980.200 ;
        RECT 4.000 976.120 1743.600 977.520 ;
        RECT 4.000 969.360 1744.010 976.120 ;
        RECT 4.400 967.960 1744.010 969.360 ;
        RECT 4.000 956.440 1744.010 967.960 ;
        RECT 4.400 955.040 1744.010 956.440 ;
        RECT 4.000 949.640 1744.010 955.040 ;
        RECT 4.000 948.240 1743.600 949.640 ;
        RECT 4.000 943.520 1744.010 948.240 ;
        RECT 4.400 942.120 1744.010 943.520 ;
        RECT 4.000 930.600 1744.010 942.120 ;
        RECT 4.400 929.200 1744.010 930.600 ;
        RECT 4.000 921.080 1744.010 929.200 ;
        RECT 4.000 919.680 1743.600 921.080 ;
        RECT 4.000 917.680 1744.010 919.680 ;
        RECT 4.400 916.280 1744.010 917.680 ;
        RECT 4.000 904.760 1744.010 916.280 ;
        RECT 4.400 903.360 1744.010 904.760 ;
        RECT 4.000 892.520 1744.010 903.360 ;
        RECT 4.000 891.840 1743.600 892.520 ;
        RECT 4.400 891.120 1743.600 891.840 ;
        RECT 4.400 890.440 1744.010 891.120 ;
        RECT 4.000 879.600 1744.010 890.440 ;
        RECT 4.400 878.200 1744.010 879.600 ;
        RECT 4.000 866.680 1744.010 878.200 ;
        RECT 4.400 865.280 1744.010 866.680 ;
        RECT 4.000 864.640 1744.010 865.280 ;
        RECT 4.000 863.240 1743.600 864.640 ;
        RECT 4.000 853.760 1744.010 863.240 ;
        RECT 4.400 852.360 1744.010 853.760 ;
        RECT 4.000 840.840 1744.010 852.360 ;
        RECT 4.400 839.440 1744.010 840.840 ;
        RECT 4.000 836.080 1744.010 839.440 ;
        RECT 4.000 834.680 1743.600 836.080 ;
        RECT 4.000 827.920 1744.010 834.680 ;
        RECT 4.400 826.520 1744.010 827.920 ;
        RECT 4.000 815.000 1744.010 826.520 ;
        RECT 4.400 813.600 1744.010 815.000 ;
        RECT 4.000 807.520 1744.010 813.600 ;
        RECT 4.000 806.120 1743.600 807.520 ;
        RECT 4.000 802.080 1744.010 806.120 ;
        RECT 4.400 800.680 1744.010 802.080 ;
        RECT 4.000 789.160 1744.010 800.680 ;
        RECT 4.400 787.760 1744.010 789.160 ;
        RECT 4.000 779.640 1744.010 787.760 ;
        RECT 4.000 778.240 1743.600 779.640 ;
        RECT 4.000 776.920 1744.010 778.240 ;
        RECT 4.400 775.520 1744.010 776.920 ;
        RECT 4.000 764.000 1744.010 775.520 ;
        RECT 4.400 762.600 1744.010 764.000 ;
        RECT 4.000 751.080 1744.010 762.600 ;
        RECT 4.400 749.680 1743.600 751.080 ;
        RECT 4.000 738.160 1744.010 749.680 ;
        RECT 4.400 736.760 1744.010 738.160 ;
        RECT 4.000 725.240 1744.010 736.760 ;
        RECT 4.400 723.840 1744.010 725.240 ;
        RECT 4.000 722.520 1744.010 723.840 ;
        RECT 4.000 721.120 1743.600 722.520 ;
        RECT 4.000 712.320 1744.010 721.120 ;
        RECT 4.400 710.920 1744.010 712.320 ;
        RECT 4.000 699.400 1744.010 710.920 ;
        RECT 4.400 698.000 1744.010 699.400 ;
        RECT 4.000 694.640 1744.010 698.000 ;
        RECT 4.000 693.240 1743.600 694.640 ;
        RECT 4.000 687.160 1744.010 693.240 ;
        RECT 4.400 685.760 1744.010 687.160 ;
        RECT 4.000 674.240 1744.010 685.760 ;
        RECT 4.400 672.840 1744.010 674.240 ;
        RECT 4.000 666.080 1744.010 672.840 ;
        RECT 4.000 664.680 1743.600 666.080 ;
        RECT 4.000 661.320 1744.010 664.680 ;
        RECT 4.400 659.920 1744.010 661.320 ;
        RECT 4.000 648.400 1744.010 659.920 ;
        RECT 4.400 647.000 1744.010 648.400 ;
        RECT 4.000 637.520 1744.010 647.000 ;
        RECT 4.000 636.120 1743.600 637.520 ;
        RECT 4.000 635.480 1744.010 636.120 ;
        RECT 4.400 634.080 1744.010 635.480 ;
        RECT 4.000 622.560 1744.010 634.080 ;
        RECT 4.400 621.160 1744.010 622.560 ;
        RECT 4.000 609.640 1744.010 621.160 ;
        RECT 4.400 608.240 1743.600 609.640 ;
        RECT 4.000 596.720 1744.010 608.240 ;
        RECT 4.400 595.320 1744.010 596.720 ;
        RECT 4.000 584.480 1744.010 595.320 ;
        RECT 4.400 583.080 1744.010 584.480 ;
        RECT 4.000 581.080 1744.010 583.080 ;
        RECT 4.000 579.680 1743.600 581.080 ;
        RECT 4.000 571.560 1744.010 579.680 ;
        RECT 4.400 570.160 1744.010 571.560 ;
        RECT 4.000 558.640 1744.010 570.160 ;
        RECT 4.400 557.240 1744.010 558.640 ;
        RECT 4.000 552.520 1744.010 557.240 ;
        RECT 4.000 551.120 1743.600 552.520 ;
        RECT 4.000 545.720 1744.010 551.120 ;
        RECT 4.400 544.320 1744.010 545.720 ;
        RECT 4.000 532.800 1744.010 544.320 ;
        RECT 4.400 531.400 1744.010 532.800 ;
        RECT 4.000 524.640 1744.010 531.400 ;
        RECT 4.000 523.240 1743.600 524.640 ;
        RECT 4.000 519.880 1744.010 523.240 ;
        RECT 4.400 518.480 1744.010 519.880 ;
        RECT 4.000 506.960 1744.010 518.480 ;
        RECT 4.400 505.560 1744.010 506.960 ;
        RECT 4.000 496.080 1744.010 505.560 ;
        RECT 4.000 494.680 1743.600 496.080 ;
        RECT 4.000 494.040 1744.010 494.680 ;
        RECT 4.400 492.640 1744.010 494.040 ;
        RECT 4.000 481.800 1744.010 492.640 ;
        RECT 4.400 480.400 1744.010 481.800 ;
        RECT 4.000 468.880 1744.010 480.400 ;
        RECT 4.400 467.520 1744.010 468.880 ;
        RECT 4.400 467.480 1743.600 467.520 ;
        RECT 4.000 466.120 1743.600 467.480 ;
        RECT 4.000 455.960 1744.010 466.120 ;
        RECT 4.400 454.560 1744.010 455.960 ;
        RECT 4.000 443.040 1744.010 454.560 ;
        RECT 4.400 441.640 1744.010 443.040 ;
        RECT 4.000 439.640 1744.010 441.640 ;
        RECT 4.000 438.240 1743.600 439.640 ;
        RECT 4.000 430.120 1744.010 438.240 ;
        RECT 4.400 428.720 1744.010 430.120 ;
        RECT 4.000 417.200 1744.010 428.720 ;
        RECT 4.400 415.800 1744.010 417.200 ;
        RECT 4.000 411.080 1744.010 415.800 ;
        RECT 4.000 409.680 1743.600 411.080 ;
        RECT 4.000 404.280 1744.010 409.680 ;
        RECT 4.400 402.880 1744.010 404.280 ;
        RECT 4.000 392.040 1744.010 402.880 ;
        RECT 4.400 390.640 1744.010 392.040 ;
        RECT 4.000 382.520 1744.010 390.640 ;
        RECT 4.000 381.120 1743.600 382.520 ;
        RECT 4.000 379.120 1744.010 381.120 ;
        RECT 4.400 377.720 1744.010 379.120 ;
        RECT 4.000 366.200 1744.010 377.720 ;
        RECT 4.400 364.800 1744.010 366.200 ;
        RECT 4.000 354.640 1744.010 364.800 ;
        RECT 4.000 353.280 1743.600 354.640 ;
        RECT 4.400 353.240 1743.600 353.280 ;
        RECT 4.400 351.880 1744.010 353.240 ;
        RECT 4.000 340.360 1744.010 351.880 ;
        RECT 4.400 338.960 1744.010 340.360 ;
        RECT 4.000 327.440 1744.010 338.960 ;
        RECT 4.400 326.080 1744.010 327.440 ;
        RECT 4.400 326.040 1743.600 326.080 ;
        RECT 4.000 324.680 1743.600 326.040 ;
        RECT 4.000 314.520 1744.010 324.680 ;
        RECT 4.400 313.120 1744.010 314.520 ;
        RECT 4.000 301.600 1744.010 313.120 ;
        RECT 4.400 300.200 1744.010 301.600 ;
        RECT 4.000 297.520 1744.010 300.200 ;
        RECT 4.000 296.120 1743.600 297.520 ;
        RECT 4.000 289.360 1744.010 296.120 ;
        RECT 4.400 287.960 1744.010 289.360 ;
        RECT 4.000 276.440 1744.010 287.960 ;
        RECT 4.400 275.040 1744.010 276.440 ;
        RECT 4.000 269.640 1744.010 275.040 ;
        RECT 4.000 268.240 1743.600 269.640 ;
        RECT 4.000 263.520 1744.010 268.240 ;
        RECT 4.400 262.120 1744.010 263.520 ;
        RECT 4.000 250.600 1744.010 262.120 ;
        RECT 4.400 249.200 1744.010 250.600 ;
        RECT 4.000 241.080 1744.010 249.200 ;
        RECT 4.000 239.680 1743.600 241.080 ;
        RECT 4.000 237.680 1744.010 239.680 ;
        RECT 4.400 236.280 1744.010 237.680 ;
        RECT 4.000 224.760 1744.010 236.280 ;
        RECT 4.400 223.360 1744.010 224.760 ;
        RECT 4.000 212.520 1744.010 223.360 ;
        RECT 4.000 211.840 1743.600 212.520 ;
        RECT 4.400 211.120 1743.600 211.840 ;
        RECT 4.400 210.440 1744.010 211.120 ;
        RECT 4.000 199.600 1744.010 210.440 ;
        RECT 4.400 198.200 1744.010 199.600 ;
        RECT 4.000 186.680 1744.010 198.200 ;
        RECT 4.400 185.280 1744.010 186.680 ;
        RECT 4.000 184.640 1744.010 185.280 ;
        RECT 4.000 183.240 1743.600 184.640 ;
        RECT 4.000 173.760 1744.010 183.240 ;
        RECT 4.400 172.360 1744.010 173.760 ;
        RECT 4.000 160.840 1744.010 172.360 ;
        RECT 4.400 159.440 1744.010 160.840 ;
        RECT 4.000 156.080 1744.010 159.440 ;
        RECT 4.000 154.680 1743.600 156.080 ;
        RECT 4.000 147.920 1744.010 154.680 ;
        RECT 4.400 146.520 1744.010 147.920 ;
        RECT 4.000 135.000 1744.010 146.520 ;
        RECT 4.400 133.600 1744.010 135.000 ;
        RECT 4.000 127.520 1744.010 133.600 ;
        RECT 4.000 126.120 1743.600 127.520 ;
        RECT 4.000 122.080 1744.010 126.120 ;
        RECT 4.400 120.680 1744.010 122.080 ;
        RECT 4.000 109.160 1744.010 120.680 ;
        RECT 4.400 107.760 1744.010 109.160 ;
        RECT 4.000 99.640 1744.010 107.760 ;
        RECT 4.000 98.240 1743.600 99.640 ;
        RECT 4.000 96.920 1744.010 98.240 ;
        RECT 4.400 95.520 1744.010 96.920 ;
        RECT 4.000 84.000 1744.010 95.520 ;
        RECT 4.400 82.600 1744.010 84.000 ;
        RECT 4.000 71.080 1744.010 82.600 ;
        RECT 4.400 69.680 1743.600 71.080 ;
        RECT 4.000 58.160 1744.010 69.680 ;
        RECT 4.400 56.760 1744.010 58.160 ;
        RECT 4.000 45.240 1744.010 56.760 ;
        RECT 4.400 43.840 1744.010 45.240 ;
        RECT 4.000 42.520 1744.010 43.840 ;
        RECT 4.000 41.120 1743.600 42.520 ;
        RECT 4.000 32.320 1744.010 41.120 ;
        RECT 4.400 30.920 1744.010 32.320 ;
        RECT 4.000 19.400 1744.010 30.920 ;
        RECT 4.400 18.000 1744.010 19.400 ;
        RECT 4.000 14.640 1744.010 18.000 ;
        RECT 4.000 13.240 1743.600 14.640 ;
        RECT 4.000 7.160 1744.010 13.240 ;
        RECT 4.400 6.295 1744.010 7.160 ;
      LAYER met4 ;
        RECT 4.895 10.640 1736.170 1349.360 ;
  END
END pyfive_top
END LIBRARY

